module lp_40x40_rom(
    input  [5:0] x_idx,
    input  [5:0] y_idx,
    output reg [7:0] RED,
    output reg [7:0] GRN,
    output reg [7:0] BLU);
always @ (*)
    case ({y_idx,x_idx})
        0:
        begin
            RED=8'h01;
            GRN=8'h01;
            BLU=8'h01;
        end
        1:
        begin
            RED=8'h01;
            GRN=8'h01;
            BLU=8'h01;
        end
        2:
        begin
            RED=8'h02;
            GRN=8'h02;
            BLU=8'h04;
        end
        3:
        begin
            RED=8'h02;
            GRN=8'h02;
            BLU=8'h04;
        end
        4:
        begin
            RED=8'h03;
            GRN=8'h02;
            BLU=8'h08;
        end
        5:
        begin
            RED=8'h02;
            GRN=8'h01;
            BLU=8'h07;
        end
        6:
        begin
            RED=8'h04;
            GRN=8'h03;
            BLU=8'h09;
        end
        7:
        begin
            RED=8'h05;
            GRN=8'h04;
            BLU=8'h0A;
        end
        8:
        begin
            RED=8'h07;
            GRN=8'h07;
            BLU=8'h09;
        end
        9:
        begin
            RED=8'h07;
            GRN=8'h06;
            BLU=8'h0E;
        end
        10:
        begin
            RED=8'h09;
            GRN=8'h07;
            BLU=8'h12;
        end
        11:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        12:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        13:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        14:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        15:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        16:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        17:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h13;
        end
        18:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h13;
        end
        19:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h13;
        end
        20:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h14;
        end
        21:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h13;
        end
        22:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h15;
        end
        23:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        24:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        25:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        26:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        27:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        28:
        begin
            RED=8'h07;
            GRN=8'h06;
            BLU=8'h0E;
        end
        29:
        begin
            RED=8'h08;
            GRN=8'h07;
            BLU=8'h0C;
        end
        30:
        begin
            RED=8'h06;
            GRN=8'h06;
            BLU=8'h08;
        end
        31:
        begin
            RED=8'h05;
            GRN=8'h04;
            BLU=8'h09;
        end
        32:
        begin
            RED=8'h04;
            GRN=8'h03;
            BLU=8'h09;
        end
        33:
        begin
            RED=8'h03;
            GRN=8'h02;
            BLU=8'h07;
        end
        34:
        begin
            RED=8'h02;
            GRN=8'h02;
            BLU=8'h04;
        end
        35:
        begin
            RED=8'h02;
            GRN=8'h02;
            BLU=8'h02;
        end
        36:
        begin
            RED=8'h01;
            GRN=8'h01;
            BLU=8'h01;
        end
        37:
        begin
            RED=8'h01;
            GRN=8'h01;
            BLU=8'h01;
        end
        38:
        begin
            RED=8'h01;
            GRN=8'h01;
            BLU=8'h01;
        end
        39:
        begin
            RED=8'h01;
            GRN=8'h01;
            BLU=8'h01;
        end
        64:
        begin
            RED=8'h01;
            GRN=8'h01;
            BLU=8'h01;
        end
        65:
        begin
            RED=8'h02;
            GRN=8'h02;
            BLU=8'h04;
        end
        66:
        begin
            RED=8'h02;
            GRN=8'h02;
            BLU=8'h04;
        end
        67:
        begin
            RED=8'h02;
            GRN=8'h02;
            BLU=8'h04;
        end
        68:
        begin
            RED=8'h03;
            GRN=8'h02;
            BLU=8'h08;
        end
        69:
        begin
            RED=8'h04;
            GRN=8'h03;
            BLU=8'h09;
        end
        70:
        begin
            RED=8'h05;
            GRN=8'h04;
            BLU=8'h0A;
        end
        71:
        begin
            RED=8'h07;
            GRN=8'h06;
            BLU=8'h0E;
        end
        72:
        begin
            RED=8'h08;
            GRN=8'h07;
            BLU=8'h0C;
        end
        73:
        begin
            RED=8'h09;
            GRN=8'h08;
            BLU=8'h10;
        end
        74:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        75:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        76:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h15;
        end
        77:
        begin
            RED=8'h0C;
            GRN=8'h0B;
            BLU=8'h13;
        end
        78:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h15;
        end
        79:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h13;
        end
        80:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h13;
        end
        81:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h16;
        end
        82:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h14;
        end
        83:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        84:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h14;
        end
        85:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h16;
        end
        86:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h14;
        end
        87:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h13;
        end
        88:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h13;
        end
        89:
        begin
            RED=8'h0C;
            GRN=8'h0B;
            BLU=8'h13;
        end
        90:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        91:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        92:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h0F;
        end
        93:
        begin
            RED=8'h08;
            GRN=8'h07;
            BLU=8'h0C;
        end
        94:
        begin
            RED=8'h07;
            GRN=8'h06;
            BLU=8'h0C;
        end
        95:
        begin
            RED=8'h06;
            GRN=8'h05;
            BLU=8'h0A;
        end
        96:
        begin
            RED=8'h05;
            GRN=8'h05;
            BLU=8'h07;
        end
        97:
        begin
            RED=8'h04;
            GRN=8'h03;
            BLU=8'h08;
        end
        98:
        begin
            RED=8'h03;
            GRN=8'h03;
            BLU=8'h05;
        end
        99:
        begin
            RED=8'h03;
            GRN=8'h03;
            BLU=8'h05;
        end
        100:
        begin
            RED=8'h02;
            GRN=8'h02;
            BLU=8'h02;
        end
        101:
        begin
            RED=8'h01;
            GRN=8'h01;
            BLU=8'h01;
        end
        102:
        begin
            RED=8'h01;
            GRN=8'h01;
            BLU=8'h01;
        end
        103:
        begin
            RED=8'h01;
            GRN=8'h01;
            BLU=8'h01;
        end
        128:
        begin
            RED=8'h02;
            GRN=8'h02;
            BLU=8'h04;
        end
        129:
        begin
            RED=8'h02;
            GRN=8'h02;
            BLU=8'h04;
        end
        130:
        begin
            RED=8'h03;
            GRN=8'h03;
            BLU=8'h05;
        end
        131:
        begin
            RED=8'h03;
            GRN=8'h02;
            BLU=8'h07;
        end
        132:
        begin
            RED=8'h04;
            GRN=8'h03;
            BLU=8'h09;
        end
        133:
        begin
            RED=8'h05;
            GRN=8'h04;
            BLU=8'h0A;
        end
        134:
        begin
            RED=8'h06;
            GRN=8'h05;
            BLU=8'h0D;
        end
        135:
        begin
            RED=8'h09;
            GRN=8'h08;
            BLU=8'h0E;
        end
        136:
        begin
            RED=8'h09;
            GRN=8'h08;
            BLU=8'h10;
        end
        137:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        138:
        begin
            RED=8'h0C;
            GRN=8'h0B;
            BLU=8'h13;
        end
        139:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h15;
        end
        140:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h14;
        end
        141:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h15;
        end
        142:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h14;
        end
        143:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h16;
        end
        144:
        begin
            RED=8'h11;
            GRN=8'h10;
            BLU=8'h18;
        end
        145:
        begin
            RED=8'h12;
            GRN=8'h11;
            BLU=8'h17;
        end
        146:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        147:
        begin
            RED=8'h11;
            GRN=8'h10;
            BLU=8'h16;
        end
        148:
        begin
            RED=8'h12;
            GRN=8'h11;
            BLU=8'h19;
        end
        149:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        150:
        begin
            RED=8'h11;
            GRN=8'h10;
            BLU=8'h16;
        end
        151:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h15;
        end
        152:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h15;
        end
        153:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h14;
        end
        154:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h16;
        end
        155:
        begin
            RED=8'h0C;
            GRN=8'h0B;
            BLU=8'h13;
        end
        156:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        157:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        158:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h0F;
        end
        159:
        begin
            RED=8'h08;
            GRN=8'h07;
            BLU=8'h0C;
        end
        160:
        begin
            RED=8'h07;
            GRN=8'h06;
            BLU=8'h0B;
        end
        161:
        begin
            RED=8'h05;
            GRN=8'h04;
            BLU=8'h09;
        end
        162:
        begin
            RED=8'h04;
            GRN=8'h03;
            BLU=8'h09;
        end
        163:
        begin
            RED=8'h03;
            GRN=8'h03;
            BLU=8'h05;
        end
        164:
        begin
            RED=8'h02;
            GRN=8'h02;
            BLU=8'h04;
        end
        165:
        begin
            RED=8'h01;
            GRN=8'h01;
            BLU=8'h01;
        end
        166:
        begin
            RED=8'h01;
            GRN=8'h01;
            BLU=8'h01;
        end
        167:
        begin
            RED=8'h01;
            GRN=8'h01;
            BLU=8'h01;
        end
        192:
        begin
            RED=8'h02;
            GRN=8'h02;
            BLU=8'h04;
        end
        193:
        begin
            RED=8'h03;
            GRN=8'h03;
            BLU=8'h05;
        end
        194:
        begin
            RED=8'h03;
            GRN=8'h02;
            BLU=8'h08;
        end
        195:
        begin
            RED=8'h04;
            GRN=8'h03;
            BLU=8'h09;
        end
        196:
        begin
            RED=8'h05;
            GRN=8'h04;
            BLU=8'h0A;
        end
        197:
        begin
            RED=8'h06;
            GRN=8'h05;
            BLU=8'h0D;
        end
        198:
        begin
            RED=8'h08;
            GRN=8'h07;
            BLU=8'h0F;
        end
        199:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        200:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        201:
        begin
            RED=8'h0C;
            GRN=8'h0B;
            BLU=8'h13;
        end
        202:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h16;
        end
        203:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h14;
        end
        204:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h15;
        end
        205:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        206:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        207:
        begin
            RED=8'h11;
            GRN=8'h10;
            BLU=8'h18;
        end
        208:
        begin
            RED=8'h12;
            GRN=8'h11;
            BLU=8'h17;
        end
        209:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h1A;
        end
        210:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h18;
        end
        211:
        begin
            RED=8'h13;
            GRN=8'h13;
            BLU=8'h15;
        end
        212:
        begin
            RED=8'h17;
            GRN=8'h16;
            BLU=8'h1C;
        end
        213:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h15;
        end
        214:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h18;
        end
        215:
        begin
            RED=8'h11;
            GRN=8'h10;
            BLU=8'h18;
        end
        216:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        217:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        218:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h14;
        end
        219:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h14;
        end
        220:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        221:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        222:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        223:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        224:
        begin
            RED=8'h08;
            GRN=8'h07;
            BLU=8'h0C;
        end
        225:
        begin
            RED=8'h05;
            GRN=8'h06;
            BLU=8'h0A;
        end
        226:
        begin
            RED=8'h04;
            GRN=8'h03;
            BLU=8'h0B;
        end
        227:
        begin
            RED=8'h02;
            GRN=8'h01;
            BLU=8'h07;
        end
        228:
        begin
            RED=8'h02;
            GRN=8'h02;
            BLU=8'h04;
        end
        229:
        begin
            RED=8'h02;
            GRN=8'h02;
            BLU=8'h04;
        end
        230:
        begin
            RED=8'h01;
            GRN=8'h01;
            BLU=8'h03;
        end
        231:
        begin
            RED=8'h01;
            GRN=8'h01;
            BLU=8'h01;
        end
        256:
        begin
            RED=8'h03;
            GRN=8'h03;
            BLU=8'h05;
        end
        257:
        begin
            RED=8'h03;
            GRN=8'h02;
            BLU=8'h08;
        end
        258:
        begin
            RED=8'h04;
            GRN=8'h03;
            BLU=8'h09;
        end
        259:
        begin
            RED=8'h04;
            GRN=8'h03;
            BLU=8'h09;
        end
        260:
        begin
            RED=8'h05;
            GRN=8'h04;
            BLU=8'h0C;
        end
        261:
        begin
            RED=8'h08;
            GRN=8'h07;
            BLU=8'h0F;
        end
        262:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        263:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        264:
        begin
            RED=8'h0C;
            GRN=8'h0B;
            BLU=8'h13;
        end
        265:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h13;
        end
        266:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        267:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h15;
        end
        268:
        begin
            RED=8'h12;
            GRN=8'h11;
            BLU=8'h19;
        end
        269:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h1A;
        end
        270:
        begin
            RED=8'h12;
            GRN=8'h11;
            BLU=8'h19;
        end
        271:
        begin
            RED=8'h14;
            GRN=8'h13;
            BLU=8'h1B;
        end
        272:
        begin
            RED=8'h14;
            GRN=8'h13;
            BLU=8'h19;
        end
        273:
        begin
            RED=8'h27;
            GRN=8'h1D;
            BLU=8'h1B;
        end
        274:
        begin
            RED=8'h43;
            GRN=8'h30;
            BLU=8'h22;
        end
        275:
        begin
            RED=8'h52;
            GRN=8'h38;
            BLU=8'h29;
        end
        276:
        begin
            RED=8'h5F;
            GRN=8'h3E;
            BLU=8'h2D;
        end
        277:
        begin
            RED=8'h4B;
            GRN=8'h37;
            BLU=8'h2C;
        end
        278:
        begin
            RED=8'h3C;
            GRN=8'h2E;
            BLU=8'h23;
        end
        279:
        begin
            RED=8'h11;
            GRN=8'h11;
            BLU=8'h1B;
        end
        280:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h18;
        end
        281:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h18;
        end
        282:
        begin
            RED=8'h11;
            GRN=8'h10;
            BLU=8'h16;
        end
        283:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        284:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h15;
        end
        285:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        286:
        begin
            RED=8'h0C;
            GRN=8'h0B;
            BLU=8'h13;
        end
        287:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        288:
        begin
            RED=8'h09;
            GRN=8'h08;
            BLU=8'h0D;
        end
        289:
        begin
            RED=8'h07;
            GRN=8'h07;
            BLU=8'h09;
        end
        290:
        begin
            RED=8'h06;
            GRN=8'h07;
            BLU=8'h0C;
        end
        291:
        begin
            RED=8'h04;
            GRN=8'h03;
            BLU=8'h09;
        end
        292:
        begin
            RED=8'h03;
            GRN=8'h03;
            BLU=8'h05;
        end
        293:
        begin
            RED=8'h02;
            GRN=8'h02;
            BLU=8'h04;
        end
        294:
        begin
            RED=8'h02;
            GRN=8'h02;
            BLU=8'h04;
        end
        295:
        begin
            RED=8'h01;
            GRN=8'h01;
            BLU=8'h01;
        end
        320:
        begin
            RED=8'h03;
            GRN=8'h03;
            BLU=8'h03;
        end
        321:
        begin
            RED=8'h03;
            GRN=8'h02;
            BLU=8'h08;
        end
        322:
        begin
            RED=8'h04;
            GRN=8'h03;
            BLU=8'h09;
        end
        323:
        begin
            RED=8'h06;
            GRN=8'h05;
            BLU=8'h0B;
        end
        324:
        begin
            RED=8'h06;
            GRN=8'h05;
            BLU=8'h0D;
        end
        325:
        begin
            RED=8'h09;
            GRN=8'h08;
            BLU=8'h10;
        end
        326:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        327:
        begin
            RED=8'h0C;
            GRN=8'h0B;
            BLU=8'h13;
        end
        328:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h13;
        end
        329:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h14;
        end
        330:
        begin
            RED=8'h11;
            GRN=8'h10;
            BLU=8'h16;
        end
        331:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h1A;
        end
        332:
        begin
            RED=8'h14;
            GRN=8'h13;
            BLU=8'h1B;
        end
        333:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h1A;
        end
        334:
        begin
            RED=8'h14;
            GRN=8'h13;
            BLU=8'h1B;
        end
        335:
        begin
            RED=8'h15;
            GRN=8'h14;
            BLU=8'h1C;
        end
        336:
        begin
            RED=8'h3D;
            GRN=8'h29;
            BLU=8'h20;
        end
        337:
        begin
            RED=8'h73;
            GRN=8'h53;
            BLU=8'h44;
        end
        338:
        begin
            RED=8'hA8;
            GRN=8'h7F;
            BLU=8'h69;
        end
        339:
        begin
            RED=8'hA5;
            GRN=8'h78;
            BLU=8'h61;
        end
        340:
        begin
            RED=8'hB8;
            GRN=8'h86;
            BLU=8'h6D;
        end
        341:
        begin
            RED=8'hAC;
            GRN=8'h7E;
            BLU=8'h67;
        end
        342:
        begin
            RED=8'h88;
            GRN=8'h65;
            BLU=8'h51;
        end
        343:
        begin
            RED=8'h78;
            GRN=8'h57;
            BLU=8'h46;
        end
        344:
        begin
            RED=8'h32;
            GRN=8'h2A;
            BLU=8'h27;
        end
        345:
        begin
            RED=8'h12;
            GRN=8'h11;
            BLU=8'h17;
        end
        346:
        begin
            RED=8'h12;
            GRN=8'h11;
            BLU=8'h17;
        end
        347:
        begin
            RED=8'h12;
            GRN=8'h11;
            BLU=8'h17;
        end
        348:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h15;
        end
        349:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h13;
        end
        350:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        351:
        begin
            RED=8'h0C;
            GRN=8'h0B;
            BLU=8'h13;
        end
        352:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        353:
        begin
            RED=8'h09;
            GRN=8'h08;
            BLU=8'h0D;
        end
        354:
        begin
            RED=8'h08;
            GRN=8'h07;
            BLU=8'h0F;
        end
        355:
        begin
            RED=8'h05;
            GRN=8'h04;
            BLU=8'h09;
        end
        356:
        begin
            RED=8'h04;
            GRN=8'h03;
            BLU=8'h09;
        end
        357:
        begin
            RED=8'h03;
            GRN=8'h03;
            BLU=8'h05;
        end
        358:
        begin
            RED=8'h02;
            GRN=8'h02;
            BLU=8'h04;
        end
        359:
        begin
            RED=8'h02;
            GRN=8'h02;
            BLU=8'h02;
        end
        384:
        begin
            RED=8'h03;
            GRN=8'h03;
            BLU=8'h03;
        end
        385:
        begin
            RED=8'h04;
            GRN=8'h03;
            BLU=8'h09;
        end
        386:
        begin
            RED=8'h05;
            GRN=8'h04;
            BLU=8'h0A;
        end
        387:
        begin
            RED=8'h07;
            GRN=8'h06;
            BLU=8'h0E;
        end
        388:
        begin
            RED=8'h09;
            GRN=8'h08;
            BLU=8'h10;
        end
        389:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        390:
        begin
            RED=8'h0C;
            GRN=8'h0B;
            BLU=8'h13;
        end
        391:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h13;
        end
        392:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        393:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h16;
        end
        394:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h1A;
        end
        395:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h1A;
        end
        396:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h1A;
        end
        397:
        begin
            RED=8'h15;
            GRN=8'h14;
            BLU=8'h1C;
        end
        398:
        begin
            RED=8'h15;
            GRN=8'h12;
            BLU=8'h19;
        end
        399:
        begin
            RED=8'h37;
            GRN=8'h25;
            BLU=8'h1B;
        end
        400:
        begin
            RED=8'hBC;
            GRN=8'h85;
            BLU=8'h67;
        end
        401:
        begin
            RED=8'hCF;
            GRN=8'h93;
            BLU=8'h77;
        end
        402:
        begin
            RED=8'hDB;
            GRN=8'h9A;
            BLU=8'h7E;
        end
        403:
        begin
            RED=8'hDF;
            GRN=8'h9E;
            BLU=8'h80;
        end
        404:
        begin
            RED=8'hE5;
            GRN=8'hA2;
            BLU=8'h85;
        end
        405:
        begin
            RED=8'hE6;
            GRN=8'hA4;
            BLU=8'h84;
        end
        406:
        begin
            RED=8'hD9;
            GRN=8'h98;
            BLU=8'h7A;
        end
        407:
        begin
            RED=8'hCF;
            GRN=8'h96;
            BLU=8'h79;
        end
        408:
        begin
            RED=8'hA1;
            GRN=8'h71;
            BLU=8'h5A;
        end
        409:
        begin
            RED=8'h2E;
            GRN=8'h29;
            BLU=8'h23;
        end
        410:
        begin
            RED=8'h12;
            GRN=8'h11;
            BLU=8'h19;
        end
        411:
        begin
            RED=8'h14;
            GRN=8'h13;
            BLU=8'h1B;
        end
        412:
        begin
            RED=8'h12;
            GRN=8'h11;
            BLU=8'h19;
        end
        413:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h15;
        end
        414:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h15;
        end
        415:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h15;
        end
        416:
        begin
            RED=8'h0C;
            GRN=8'h0B;
            BLU=8'h13;
        end
        417:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        418:
        begin
            RED=8'h07;
            GRN=8'h07;
            BLU=8'h09;
        end
        419:
        begin
            RED=8'h06;
            GRN=8'h05;
            BLU=8'h0D;
        end
        420:
        begin
            RED=8'h04;
            GRN=8'h04;
            BLU=8'h06;
        end
        421:
        begin
            RED=8'h03;
            GRN=8'h02;
            BLU=8'h08;
        end
        422:
        begin
            RED=8'h03;
            GRN=8'h03;
            BLU=8'h05;
        end
        423:
        begin
            RED=8'h02;
            GRN=8'h02;
            BLU=8'h04;
        end
        448:
        begin
            RED=8'h04;
            GRN=8'h03;
            BLU=8'h09;
        end
        449:
        begin
            RED=8'h04;
            GRN=8'h03;
            BLU=8'h09;
        end
        450:
        begin
            RED=8'h06;
            GRN=8'h05;
            BLU=8'h0D;
        end
        451:
        begin
            RED=8'h09;
            GRN=8'h08;
            BLU=8'h10;
        end
        452:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        453:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        454:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h15;
        end
        455:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h16;
        end
        456:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        457:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h1A;
        end
        458:
        begin
            RED=8'h14;
            GRN=8'h13;
            BLU=8'h1B;
        end
        459:
        begin
            RED=8'h14;
            GRN=8'h13;
            BLU=8'h1B;
        end
        460:
        begin
            RED=8'h14;
            GRN=8'h13;
            BLU=8'h1B;
        end
        461:
        begin
            RED=8'h16;
            GRN=8'h15;
            BLU=8'h1D;
        end
        462:
        begin
            RED=8'h39;
            GRN=8'h28;
            BLU=8'h20;
        end
        463:
        begin
            RED=8'hBF;
            GRN=8'h87;
            BLU=8'h6E;
        end
        464:
        begin
            RED=8'hCE;
            GRN=8'h8E;
            BLU=8'h72;
        end
        465:
        begin
            RED=8'hE0;
            GRN=8'h96;
            BLU=8'h79;
        end
        466:
        begin
            RED=8'hE6;
            GRN=8'h9F;
            BLU=8'h83;
        end
        467:
        begin
            RED=8'hEB;
            GRN=8'hA4;
            BLU=8'h88;
        end
        468:
        begin
            RED=8'hF5;
            GRN=8'hAB;
            BLU=8'h8E;
        end
        469:
        begin
            RED=8'hEB;
            GRN=8'hA4;
            BLU=8'h88;
        end
        470:
        begin
            RED=8'hE8;
            GRN=8'hA1;
            BLU=8'h83;
        end
        471:
        begin
            RED=8'hDE;
            GRN=8'h9C;
            BLU=8'h7C;
        end
        472:
        begin
            RED=8'hCE;
            GRN=8'h93;
            BLU=8'h73;
        end
        473:
        begin
            RED=8'hB0;
            GRN=8'h81;
            BLU=8'h67;
        end
        474:
        begin
            RED=8'h31;
            GRN=8'h2D;
            BLU=8'h2E;
        end
        475:
        begin
            RED=8'h14;
            GRN=8'h13;
            BLU=8'h1B;
        end
        476:
        begin
            RED=8'h12;
            GRN=8'h11;
            BLU=8'h17;
        end
        477:
        begin
            RED=8'h11;
            GRN=8'h10;
            BLU=8'h18;
        end
        478:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        479:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h15;
        end
        480:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        481:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        482:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        483:
        begin
            RED=8'h09;
            GRN=8'h08;
            BLU=8'h0E;
        end
        484:
        begin
            RED=8'h07;
            GRN=8'h07;
            BLU=8'h09;
        end
        485:
        begin
            RED=8'h03;
            GRN=8'h02;
            BLU=8'h08;
        end
        486:
        begin
            RED=8'h03;
            GRN=8'h02;
            BLU=8'h0A;
        end
        487:
        begin
            RED=8'h02;
            GRN=8'h02;
            BLU=8'h04;
        end
        512:
        begin
            RED=8'h04;
            GRN=8'h03;
            BLU=8'h09;
        end
        513:
        begin
            RED=8'h05;
            GRN=8'h04;
            BLU=8'h0A;
        end
        514:
        begin
            RED=8'h08;
            GRN=8'h07;
            BLU=8'h0F;
        end
        515:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        516:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        517:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        518:
        begin
            RED=8'h11;
            GRN=8'h10;
            BLU=8'h18;
        end
        519:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        520:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h1A;
        end
        521:
        begin
            RED=8'h14;
            GRN=8'h13;
            BLU=8'h1B;
        end
        522:
        begin
            RED=8'h15;
            GRN=8'h13;
            BLU=8'h1E;
        end
        523:
        begin
            RED=8'h15;
            GRN=8'h14;
            BLU=8'h1C;
        end
        524:
        begin
            RED=8'h15;
            GRN=8'h14;
            BLU=8'h1A;
        end
        525:
        begin
            RED=8'h36;
            GRN=8'h32;
            BLU=8'h29;
        end
        526:
        begin
            RED=8'h59;
            GRN=8'h41;
            BLU=8'h35;
        end
        527:
        begin
            RED=8'hCB;
            GRN=8'h90;
            BLU=8'h72;
        end
        528:
        begin
            RED=8'hDB;
            GRN=8'h96;
            BLU=8'h79;
        end
        529:
        begin
            RED=8'hE3;
            GRN=8'h9C;
            BLU=8'h7E;
        end
        530:
        begin
            RED=8'hEC;
            GRN=8'hA7;
            BLU=8'h8A;
        end
        531:
        begin
            RED=8'hF0;
            GRN=8'hA6;
            BLU=8'h89;
        end
        532:
        begin
            RED=8'hF3;
            GRN=8'hB0;
            BLU=8'h95;
        end
        533:
        begin
            RED=8'hF0;
            GRN=8'hAE;
            BLU=8'h8E;
        end
        534:
        begin
            RED=8'hEC;
            GRN=8'hA1;
            BLU=8'h84;
        end
        535:
        begin
            RED=8'hE6;
            GRN=8'h9D;
            BLU=8'h7D;
        end
        536:
        begin
            RED=8'hD6;
            GRN=8'h96;
            BLU=8'h7A;
        end
        537:
        begin
            RED=8'hCB;
            GRN=8'h94;
            BLU=8'h75;
        end
        538:
        begin
            RED=8'h3D;
            GRN=8'h26;
            BLU=8'h18;
        end
        539:
        begin
            RED=8'h17;
            GRN=8'h16;
            BLU=8'h1C;
        end
        540:
        begin
            RED=8'h14;
            GRN=8'h13;
            BLU=8'h1B;
        end
        541:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h1A;
        end
        542:
        begin
            RED=8'h12;
            GRN=8'h11;
            BLU=8'h19;
        end
        543:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        544:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h13;
        end
        545:
        begin
            RED=8'h0C;
            GRN=8'h0B;
            BLU=8'h13;
        end
        546:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        547:
        begin
            RED=8'h09;
            GRN=8'h08;
            BLU=8'h10;
        end
        548:
        begin
            RED=8'h06;
            GRN=8'h05;
            BLU=8'h0D;
        end
        549:
        begin
            RED=8'h05;
            GRN=8'h05;
            BLU=8'h07;
        end
        550:
        begin
            RED=8'h04;
            GRN=8'h03;
            BLU=8'h09;
        end
        551:
        begin
            RED=8'h03;
            GRN=8'h02;
            BLU=8'h07;
        end
        576:
        begin
            RED=8'h05;
            GRN=8'h04;
            BLU=8'h0A;
        end
        577:
        begin
            RED=8'h06;
            GRN=8'h05;
            BLU=8'h0B;
        end
        578:
        begin
            RED=8'h09;
            GRN=8'h08;
            BLU=8'h10;
        end
        579:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        580:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h15;
        end
        581:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h13;
        end
        582:
        begin
            RED=8'h12;
            GRN=8'h11;
            BLU=8'h19;
        end
        583:
        begin
            RED=8'h12;
            GRN=8'h13;
            BLU=8'h18;
        end
        584:
        begin
            RED=8'h13;
            GRN=8'h13;
            BLU=8'h1B;
        end
        585:
        begin
            RED=8'h15;
            GRN=8'h14;
            BLU=8'h1C;
        end
        586:
        begin
            RED=8'h16;
            GRN=8'h14;
            BLU=8'h21;
        end
        587:
        begin
            RED=8'h18;
            GRN=8'h16;
            BLU=8'h21;
        end
        588:
        begin
            RED=8'h15;
            GRN=8'h13;
            BLU=8'h21;
        end
        589:
        begin
            RED=8'h52;
            GRN=8'h48;
            BLU=8'h3F;
        end
        590:
        begin
            RED=8'hAE;
            GRN=8'h84;
            BLU=8'h6C;
        end
        591:
        begin
            RED=8'hC9;
            GRN=8'h8E;
            BLU=8'h70;
        end
        592:
        begin
            RED=8'hE2;
            GRN=8'hA1;
            BLU=8'h83;
        end
        593:
        begin
            RED=8'hE6;
            GRN=8'hA5;
            BLU=8'h89;
        end
        594:
        begin
            RED=8'hE8;
            GRN=8'hA7;
            BLU=8'h8B;
        end
        595:
        begin
            RED=8'hEF;
            GRN=8'hA8;
            BLU=8'h8C;
        end
        596:
        begin
            RED=8'hEB;
            GRN=8'hAA;
            BLU=8'h8E;
        end
        597:
        begin
            RED=8'hF5;
            GRN=8'hB0;
            BLU=8'h91;
        end
        598:
        begin
            RED=8'hE6;
            GRN=8'hA1;
            BLU=8'h82;
        end
        599:
        begin
            RED=8'hE2;
            GRN=8'h9F;
            BLU=8'h82;
        end
        600:
        begin
            RED=8'hDB;
            GRN=8'h99;
            BLU=8'h79;
        end
        601:
        begin
            RED=8'hD7;
            GRN=8'h9A;
            BLU=8'h7D;
        end
        602:
        begin
            RED=8'hB6;
            GRN=8'h8A;
            BLU=8'h6F;
        end
        603:
        begin
            RED=8'h2C;
            GRN=8'h2C;
            BLU=8'h2E;
        end
        604:
        begin
            RED=8'h14;
            GRN=8'h13;
            BLU=8'h1B;
        end
        605:
        begin
            RED=8'h14;
            GRN=8'h13;
            BLU=8'h1B;
        end
        606:
        begin
            RED=8'h12;
            GRN=8'h11;
            BLU=8'h19;
        end
        607:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        608:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h14;
        end
        609:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        610:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        611:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        612:
        begin
            RED=8'h08;
            GRN=8'h08;
            BLU=8'h08;
        end
        613:
        begin
            RED=8'h05;
            GRN=8'h04;
            BLU=8'h0A;
        end
        614:
        begin
            RED=8'h04;
            GRN=8'h03;
            BLU=8'h09;
        end
        615:
        begin
            RED=8'h03;
            GRN=8'h02;
            BLU=8'h07;
        end
        640:
        begin
            RED=8'h06;
            GRN=8'h05;
            BLU=8'h0B;
        end
        641:
        begin
            RED=8'h07;
            GRN=8'h06;
            BLU=8'h0E;
        end
        642:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        643:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        644:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h14;
        end
        645:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        646:
        begin
            RED=8'h13;
            GRN=8'h11;
            BLU=8'h1C;
        end
        647:
        begin
            RED=8'h14;
            GRN=8'h13;
            BLU=8'h1B;
        end
        648:
        begin
            RED=8'h15;
            GRN=8'h14;
            BLU=8'h1A;
        end
        649:
        begin
            RED=8'h17;
            GRN=8'h15;
            BLU=8'h20;
        end
        650:
        begin
            RED=8'h18;
            GRN=8'h16;
            BLU=8'h21;
        end
        651:
        begin
            RED=8'h19;
            GRN=8'h17;
            BLU=8'h24;
        end
        652:
        begin
            RED=8'h28;
            GRN=8'h27;
            BLU=8'h2D;
        end
        653:
        begin
            RED=8'h60;
            GRN=8'h4A;
            BLU=8'h3D;
        end
        654:
        begin
            RED=8'hC6;
            GRN=8'h94;
            BLU=8'h79;
        end
        655:
        begin
            RED=8'hC8;
            GRN=8'h8B;
            BLU=8'h6E;
        end
        656:
        begin
            RED=8'hE1;
            GRN=8'hA0;
            BLU=8'h84;
        end
        657:
        begin
            RED=8'hE8;
            GRN=8'hA3;
            BLU=8'h86;
        end
        658:
        begin
            RED=8'hEE;
            GRN=8'hA7;
            BLU=8'h89;
        end
        659:
        begin
            RED=8'hF3;
            GRN=8'hAB;
            BLU=8'h92;
        end
        660:
        begin
            RED=8'hEF;
            GRN=8'hA7;
            BLU=8'h8E;
        end
        661:
        begin
            RED=8'hF5;
            GRN=8'hB0;
            BLU=8'h93;
        end
        662:
        begin
            RED=8'hEC;
            GRN=8'hA2;
            BLU=8'h85;
        end
        663:
        begin
            RED=8'hEC;
            GRN=8'hA7;
            BLU=8'h8A;
        end
        664:
        begin
            RED=8'hDE;
            GRN=8'h9C;
            BLU=8'h7C;
        end
        665:
        begin
            RED=8'hD3;
            GRN=8'h96;
            BLU=8'h79;
        end
        666:
        begin
            RED=8'hC2;
            GRN=8'h8A;
            BLU=8'h6F;
        end
        667:
        begin
            RED=8'h58;
            GRN=8'h4F;
            BLU=8'h48;
        end
        668:
        begin
            RED=8'h16;
            GRN=8'h15;
            BLU=8'h1D;
        end
        669:
        begin
            RED=8'h16;
            GRN=8'h15;
            BLU=8'h1B;
        end
        670:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h1A;
        end
        671:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h1A;
        end
        672:
        begin
            RED=8'h11;
            GRN=8'h10;
            BLU=8'h18;
        end
        673:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h14;
        end
        674:
        begin
            RED=8'h0C;
            GRN=8'h0B;
            BLU=8'h13;
        end
        675:
        begin
            RED=8'h0C;
            GRN=8'h0B;
            BLU=8'h13;
        end
        676:
        begin
            RED=8'h09;
            GRN=8'h08;
            BLU=8'h10;
        end
        677:
        begin
            RED=8'h06;
            GRN=8'h05;
            BLU=8'h0B;
        end
        678:
        begin
            RED=8'h05;
            GRN=8'h04;
            BLU=8'h0A;
        end
        679:
        begin
            RED=8'h04;
            GRN=8'h03;
            BLU=8'h09;
        end
        704:
        begin
            RED=8'h06;
            GRN=8'h05;
            BLU=8'h0D;
        end
        705:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        706:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        707:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        708:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h16;
        end
        709:
        begin
            RED=8'h11;
            GRN=8'h10;
            BLU=8'h18;
        end
        710:
        begin
            RED=8'h12;
            GRN=8'h12;
            BLU=8'h1C;
        end
        711:
        begin
            RED=8'h16;
            GRN=8'h14;
            BLU=8'h21;
        end
        712:
        begin
            RED=8'h17;
            GRN=8'h15;
            BLU=8'h23;
        end
        713:
        begin
            RED=8'h18;
            GRN=8'h16;
            BLU=8'h24;
        end
        714:
        begin
            RED=8'h18;
            GRN=8'h16;
            BLU=8'h24;
        end
        715:
        begin
            RED=8'h18;
            GRN=8'h16;
            BLU=8'h24;
        end
        716:
        begin
            RED=8'h3D;
            GRN=8'h3D;
            BLU=8'h3F;
        end
        717:
        begin
            RED=8'h72;
            GRN=8'h58;
            BLU=8'h4B;
        end
        718:
        begin
            RED=8'hC3;
            GRN=8'h94;
            BLU=8'h78;
        end
        719:
        begin
            RED=8'hCD;
            GRN=8'h90;
            BLU=8'h73;
        end
        720:
        begin
            RED=8'hE8;
            GRN=8'hA7;
            BLU=8'h89;
        end
        721:
        begin
            RED=8'hE6;
            GRN=8'hA5;
            BLU=8'h87;
        end
        722:
        begin
            RED=8'hF5;
            GRN=8'hB2;
            BLU=8'h95;
        end
        723:
        begin
            RED=8'hF7;
            GRN=8'hAF;
            BLU=8'h96;
        end
        724:
        begin
            RED=8'hF4;
            GRN=8'hB1;
            BLU=8'h96;
        end
        725:
        begin
            RED=8'hF9;
            GRN=8'hB4;
            BLU=8'h97;
        end
        726:
        begin
            RED=8'hF5;
            GRN=8'hB2;
            BLU=8'h97;
        end
        727:
        begin
            RED=8'hF0;
            GRN=8'hAA;
            BLU=8'h90;
        end
        728:
        begin
            RED=8'hE1;
            GRN=8'hA4;
            BLU=8'h85;
        end
        729:
        begin
            RED=8'hD4;
            GRN=8'h99;
            BLU=8'h79;
        end
        730:
        begin
            RED=8'hC3;
            GRN=8'h8A;
            BLU=8'h6D;
        end
        731:
        begin
            RED=8'h6C;
            GRN=8'h60;
            BLU=8'h54;
        end
        732:
        begin
            RED=8'h17;
            GRN=8'h15;
            BLU=8'h20;
        end
        733:
        begin
            RED=8'h16;
            GRN=8'h14;
            BLU=8'h22;
        end
        734:
        begin
            RED=8'h15;
            GRN=8'h13;
            BLU=8'h1E;
        end
        735:
        begin
            RED=8'h14;
            GRN=8'h13;
            BLU=8'h1B;
        end
        736:
        begin
            RED=8'h12;
            GRN=8'h11;
            BLU=8'h19;
        end
        737:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h15;
        end
        738:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h15;
        end
        739:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        740:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        741:
        begin
            RED=8'h06;
            GRN=8'h05;
            BLU=8'h0D;
        end
        742:
        begin
            RED=8'h05;
            GRN=8'h04;
            BLU=8'h0A;
        end
        743:
        begin
            RED=8'h04;
            GRN=8'h03;
            BLU=8'h09;
        end
        768:
        begin
            RED=8'h08;
            GRN=8'h07;
            BLU=8'h0F;
        end
        769:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        770:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        771:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h16;
        end
        772:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h1A;
        end
        773:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h1A;
        end
        774:
        begin
            RED=8'h15;
            GRN=8'h13;
            BLU=8'h20;
        end
        775:
        begin
            RED=8'h16;
            GRN=8'h14;
            BLU=8'h21;
        end
        776:
        begin
            RED=8'h15;
            GRN=8'h13;
            BLU=8'h21;
        end
        777:
        begin
            RED=8'h17;
            GRN=8'h15;
            BLU=8'h23;
        end
        778:
        begin
            RED=8'h18;
            GRN=8'h16;
            BLU=8'h24;
        end
        779:
        begin
            RED=8'h1A;
            GRN=8'h18;
            BLU=8'h26;
        end
        780:
        begin
            RED=8'h34;
            GRN=8'h32;
            BLU=8'h33;
        end
        781:
        begin
            RED=8'h66;
            GRN=8'h4A;
            BLU=8'h3E;
        end
        782:
        begin
            RED=8'hA5;
            GRN=8'h76;
            BLU=8'h5C;
        end
        783:
        begin
            RED=8'hCD;
            GRN=8'h8F;
            BLU=8'h76;
        end
        784:
        begin
            RED=8'hEA;
            GRN=8'hB1;
            BLU=8'h96;
        end
        785:
        begin
            RED=8'hDD;
            GRN=8'hAA;
            BLU=8'h95;
        end
        786:
        begin
            RED=8'hE6;
            GRN=8'hAC;
            BLU=8'h96;
        end
        787:
        begin
            RED=8'hE9;
            GRN=8'hA5;
            BLU=8'h8E;
        end
        788:
        begin
            RED=8'hED;
            GRN=8'hAC;
            BLU=8'h90;
        end
        789:
        begin
            RED=8'hEF;
            GRN=8'hAE;
            BLU=8'h90;
        end
        790:
        begin
            RED=8'hEC;
            GRN=8'hAB;
            BLU=8'h8F;
        end
        791:
        begin
            RED=8'hE0;
            GRN=8'h9F;
            BLU=8'h89;
        end
        792:
        begin
            RED=8'hDB;
            GRN=8'hA9;
            BLU=8'h90;
        end
        793:
        begin
            RED=8'hCF;
            GRN=8'hA1;
            BLU=8'h8A;
        end
        794:
        begin
            RED=8'hB8;
            GRN=8'h87;
            BLU=8'h69;
        end
        795:
        begin
            RED=8'h71;
            GRN=8'h67;
            BLU=8'h5D;
        end
        796:
        begin
            RED=8'h17;
            GRN=8'h15;
            BLU=8'h22;
        end
        797:
        begin
            RED=8'h17;
            GRN=8'h15;
            BLU=8'h20;
        end
        798:
        begin
            RED=8'h18;
            GRN=8'h16;
            BLU=8'h21;
        end
        799:
        begin
            RED=8'h15;
            GRN=8'h14;
            BLU=8'h1C;
        end
        800:
        begin
            RED=8'h11;
            GRN=8'h10;
            BLU=8'h18;
        end
        801:
        begin
            RED=8'h11;
            GRN=8'h10;
            BLU=8'h18;
        end
        802:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        803:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h14;
        end
        804:
        begin
            RED=8'h0C;
            GRN=8'h0B;
            BLU=8'h13;
        end
        805:
        begin
            RED=8'h09;
            GRN=8'h08;
            BLU=8'h10;
        end
        806:
        begin
            RED=8'h07;
            GRN=8'h06;
            BLU=8'h0E;
        end
        807:
        begin
            RED=8'h05;
            GRN=8'h04;
            BLU=8'h09;
        end
        832:
        begin
            RED=8'h09;
            GRN=8'h08;
            BLU=8'h10;
        end
        833:
        begin
            RED=8'h0C;
            GRN=8'h0B;
            BLU=8'h13;
        end
        834:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        835:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        836:
        begin
            RED=8'h12;
            GRN=8'h10;
            BLU=8'h1B;
        end
        837:
        begin
            RED=8'h15;
            GRN=8'h13;
            BLU=8'h20;
        end
        838:
        begin
            RED=8'h16;
            GRN=8'h14;
            BLU=8'h22;
        end
        839:
        begin
            RED=8'h18;
            GRN=8'h15;
            BLU=8'h26;
        end
        840:
        begin
            RED=8'h18;
            GRN=8'h16;
            BLU=8'h24;
        end
        841:
        begin
            RED=8'h18;
            GRN=8'h15;
            BLU=8'h26;
        end
        842:
        begin
            RED=8'h19;
            GRN=8'h18;
            BLU=8'h28;
        end
        843:
        begin
            RED=8'h1B;
            GRN=8'h18;
            BLU=8'h2B;
        end
        844:
        begin
            RED=8'h4D;
            GRN=8'h46;
            BLU=8'h3C;
        end
        845:
        begin
            RED=8'h5B;
            GRN=8'h44;
            BLU=8'h32;
        end
        846:
        begin
            RED=8'hC8;
            GRN=8'h8C;
            BLU=8'h70;
        end
        847:
        begin
            RED=8'hBF;
            GRN=8'h86;
            BLU=8'h72;
        end
        848:
        begin
            RED=8'h8B;
            GRN=8'h5C;
            BLU=8'h48;
        end
        849:
        begin
            RED=8'h94;
            GRN=8'h68;
            BLU=8'h4F;
        end
        850:
        begin
            RED=8'h85;
            GRN=8'h56;
            BLU=8'h44;
        end
        851:
        begin
            RED=8'hA9;
            GRN=8'h72;
            BLU=8'h5E;
        end
        852:
        begin
            RED=8'hC8;
            GRN=8'h83;
            BLU=8'h66;
        end
        853:
        begin
            RED=8'hD4;
            GRN=8'h91;
            BLU=8'h76;
        end
        854:
        begin
            RED=8'hC0;
            GRN=8'h7C;
            BLU=8'h65;
        end
        855:
        begin
            RED=8'h81;
            GRN=8'h54;
            BLU=8'h3F;
        end
        856:
        begin
            RED=8'h9A;
            GRN=8'h6D;
            BLU=8'h50;
        end
        857:
        begin
            RED=8'hAA;
            GRN=8'h80;
            BLU=8'h6A;
        end
        858:
        begin
            RED=8'h83;
            GRN=8'h5E;
            BLU=8'h4E;
        end
        859:
        begin
            RED=8'h5F;
            GRN=8'h50;
            BLU=8'h49;
        end
        860:
        begin
            RED=8'h19;
            GRN=8'h17;
            BLU=8'h22;
        end
        861:
        begin
            RED=8'h18;
            GRN=8'h16;
            BLU=8'h21;
        end
        862:
        begin
            RED=8'h17;
            GRN=8'h15;
            BLU=8'h20;
        end
        863:
        begin
            RED=8'h16;
            GRN=8'h14;
            BLU=8'h21;
        end
        864:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h1A;
        end
        865:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h1A;
        end
        866:
        begin
            RED=8'h11;
            GRN=8'h10;
            BLU=8'h18;
        end
        867:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h15;
        end
        868:
        begin
            RED=8'h0C;
            GRN=8'h0B;
            BLU=8'h13;
        end
        869:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        870:
        begin
            RED=8'h07;
            GRN=8'h06;
            BLU=8'h0E;
        end
        871:
        begin
            RED=8'h05;
            GRN=8'h04;
            BLU=8'h0A;
        end
        896:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        897:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        898:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h14;
        end
        899:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        900:
        begin
            RED=8'h15;
            GRN=8'h13;
            BLU=8'h20;
        end
        901:
        begin
            RED=8'h14;
            GRN=8'h12;
            BLU=8'h1F;
        end
        902:
        begin
            RED=8'h16;
            GRN=8'h14;
            BLU=8'h22;
        end
        903:
        begin
            RED=8'h18;
            GRN=8'h15;
            BLU=8'h26;
        end
        904:
        begin
            RED=8'h18;
            GRN=8'h15;
            BLU=8'h26;
        end
        905:
        begin
            RED=8'h19;
            GRN=8'h18;
            BLU=8'h2A;
        end
        906:
        begin
            RED=8'h19;
            GRN=8'h16;
            BLU=8'h29;
        end
        907:
        begin
            RED=8'h1A;
            GRN=8'h19;
            BLU=8'h2B;
        end
        908:
        begin
            RED=8'hB0;
            GRN=8'h8B;
            BLU=8'h79;
        end
        909:
        begin
            RED=8'h5B;
            GRN=8'h3B;
            BLU=8'h2E;
        end
        910:
        begin
            RED=8'hBD;
            GRN=8'h80;
            BLU=8'h64;
        end
        911:
        begin
            RED=8'h94;
            GRN=8'h66;
            BLU=8'h4F;
        end
        912:
        begin
            RED=8'hCD;
            GRN=8'h90;
            BLU=8'h74;
        end
        913:
        begin
            RED=8'h65;
            GRN=8'h3C;
            BLU=8'h28;
        end
        914:
        begin
            RED=8'h67;
            GRN=8'h3E;
            BLU=8'h2A;
        end
        915:
        begin
            RED=8'h91;
            GRN=8'h58;
            BLU=8'h3D;
        end
        916:
        begin
            RED=8'hC0;
            GRN=8'h7A;
            BLU=8'h61;
        end
        917:
        begin
            RED=8'hF9;
            GRN=8'hB7;
            BLU=8'h9D;
        end
        918:
        begin
            RED=8'hB3;
            GRN=8'h7C;
            BLU=8'h5E;
        end
        919:
        begin
            RED=8'h82;
            GRN=8'h4B;
            BLU=8'h36;
        end
        920:
        begin
            RED=8'h6B;
            GRN=8'h52;
            BLU=8'h4D;
        end
        921:
        begin
            RED=8'h45;
            GRN=8'h1B;
            BLU=8'h05;
        end
        922:
        begin
            RED=8'hA1;
            GRN=8'h78;
            BLU=8'h64;
        end
        923:
        begin
            RED=8'h57;
            GRN=8'h47;
            BLU=8'h3A;
        end
        924:
        begin
            RED=8'h1A;
            GRN=8'h18;
            BLU=8'h25;
        end
        925:
        begin
            RED=8'h18;
            GRN=8'h16;
            BLU=8'h24;
        end
        926:
        begin
            RED=8'h17;
            GRN=8'h15;
            BLU=8'h23;
        end
        927:
        begin
            RED=8'h18;
            GRN=8'h16;
            BLU=8'h23;
        end
        928:
        begin
            RED=8'h14;
            GRN=8'h12;
            BLU=8'h1D;
        end
        929:
        begin
            RED=8'h13;
            GRN=8'h11;
            BLU=8'h1C;
        end
        930:
        begin
            RED=8'h12;
            GRN=8'h11;
            BLU=8'h19;
        end
        931:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        932:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        933:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        934:
        begin
            RED=8'h08;
            GRN=8'h07;
            BLU=8'h0F;
        end
        935:
        begin
            RED=8'h06;
            GRN=8'h05;
            BLU=8'h0D;
        end
        960:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        961:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        962:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        963:
        begin
            RED=8'h13;
            GRN=8'h11;
            BLU=8'h1E;
        end
        964:
        begin
            RED=8'h15;
            GRN=8'h13;
            BLU=8'h21;
        end
        965:
        begin
            RED=8'h15;
            GRN=8'h12;
            BLU=8'h23;
        end
        966:
        begin
            RED=8'h18;
            GRN=8'h15;
            BLU=8'h26;
        end
        967:
        begin
            RED=8'h19;
            GRN=8'h16;
            BLU=8'h29;
        end
        968:
        begin
            RED=8'h18;
            GRN=8'h17;
            BLU=8'h29;
        end
        969:
        begin
            RED=8'h1A;
            GRN=8'h19;
            BLU=8'h2B;
        end
        970:
        begin
            RED=8'h19;
            GRN=8'h18;
            BLU=8'h2A;
        end
        971:
        begin
            RED=8'h1C;
            GRN=8'h1A;
            BLU=8'h2F;
        end
        972:
        begin
            RED=8'h96;
            GRN=8'h51;
            BLU=8'h41;
        end
        973:
        begin
            RED=8'h91;
            GRN=8'h66;
            BLU=8'h53;
        end
        974:
        begin
            RED=8'hC7;
            GRN=8'h87;
            BLU=8'h6C;
        end
        975:
        begin
            RED=8'hC9;
            GRN=8'h94;
            BLU=8'h75;
        end
        976:
        begin
            RED=8'hA3;
            GRN=8'h6A;
            BLU=8'h59;
        end
        977:
        begin
            RED=8'hC4;
            GRN=8'h94;
            BLU=8'h86;
        end
        978:
        begin
            RED=8'hDB;
            GRN=8'h9E;
            BLU=8'h8C;
        end
        979:
        begin
            RED=8'hDF;
            GRN=8'hAC;
            BLU=8'h8F;
        end
        980:
        begin
            RED=8'hD4;
            GRN=8'h8D;
            BLU=8'h71;
        end
        981:
        begin
            RED=8'hFA;
            GRN=8'hB7;
            BLU=8'h9C;
        end
        982:
        begin
            RED=8'hD4;
            GRN=8'h95;
            BLU=8'h74;
        end
        983:
        begin
            RED=8'hCA;
            GRN=8'h89;
            BLU=8'h6D;
        end
        984:
        begin
            RED=8'hCB;
            GRN=8'h8B;
            BLU=8'h72;
        end
        985:
        begin
            RED=8'hC5;
            GRN=8'h8F;
            BLU=8'h77;
        end
        986:
        begin
            RED=8'hD6;
            GRN=8'hA0;
            BLU=8'h7C;
        end
        987:
        begin
            RED=8'hB6;
            GRN=8'h84;
            BLU=8'h6B;
        end
        988:
        begin
            RED=8'h15;
            GRN=8'h17;
            BLU=8'h24;
        end
        989:
        begin
            RED=8'h19;
            GRN=8'h17;
            BLU=8'h25;
        end
        990:
        begin
            RED=8'h18;
            GRN=8'h16;
            BLU=8'h24;
        end
        991:
        begin
            RED=8'h17;
            GRN=8'h15;
            BLU=8'h23;
        end
        992:
        begin
            RED=8'h16;
            GRN=8'h14;
            BLU=8'h21;
        end
        993:
        begin
            RED=8'h15;
            GRN=8'h13;
            BLU=8'h1E;
        end
        994:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h1A;
        end
        995:
        begin
            RED=8'h11;
            GRN=8'h10;
            BLU=8'h18;
        end
        996:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h15;
        end
        997:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        998:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        999:
        begin
            RED=8'h07;
            GRN=8'h06;
            BLU=8'h0E;
        end
        1024:
        begin
            RED=8'h0E;
            GRN=8'h0C;
            BLU=8'h17;
        end
        1025:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h15;
        end
        1026:
        begin
            RED=8'h12;
            GRN=8'h10;
            BLU=8'h1D;
        end
        1027:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h20;
        end
        1028:
        begin
            RED=8'h16;
            GRN=8'h13;
            BLU=8'h26;
        end
        1029:
        begin
            RED=8'h16;
            GRN=8'h13;
            BLU=8'h24;
        end
        1030:
        begin
            RED=8'h18;
            GRN=8'h15;
            BLU=8'h28;
        end
        1031:
        begin
            RED=8'h1A;
            GRN=8'h17;
            BLU=8'h2C;
        end
        1032:
        begin
            RED=8'h19;
            GRN=8'h15;
            BLU=8'h2C;
        end
        1033:
        begin
            RED=8'h18;
            GRN=8'h14;
            BLU=8'h2B;
        end
        1034:
        begin
            RED=8'h1B;
            GRN=8'h17;
            BLU=8'h2E;
        end
        1035:
        begin
            RED=8'h1C;
            GRN=8'h19;
            BLU=8'h2E;
        end
        1036:
        begin
            RED=8'hC6;
            GRN=8'h88;
            BLU=8'h6F;
        end
        1037:
        begin
            RED=8'hA6;
            GRN=8'h73;
            BLU=8'h60;
        end
        1038:
        begin
            RED=8'hB9;
            GRN=8'h7E;
            BLU=8'h60;
        end
        1039:
        begin
            RED=8'hEC;
            GRN=8'hAF;
            BLU=8'h92;
        end
        1040:
        begin
            RED=8'hDE;
            GRN=8'hA5;
            BLU=8'h87;
        end
        1041:
        begin
            RED=8'hDA;
            GRN=8'h9C;
            BLU=8'h83;
        end
        1042:
        begin
            RED=8'hD7;
            GRN=8'h97;
            BLU=8'h7C;
        end
        1043:
        begin
            RED=8'hF2;
            GRN=8'hB2;
            BLU=8'h96;
        end
        1044:
        begin
            RED=8'hD6;
            GRN=8'h93;
            BLU=8'h79;
        end
        1045:
        begin
            RED=8'hFD;
            GRN=8'hB5;
            BLU=8'h9F;
        end
        1046:
        begin
            RED=8'hD2;
            GRN=8'h92;
            BLU=8'h77;
        end
        1047:
        begin
            RED=8'hE7;
            GRN=8'h9B;
            BLU=8'h83;
        end
        1048:
        begin
            RED=8'hF0;
            GRN=8'hAF;
            BLU=8'h91;
        end
        1049:
        begin
            RED=8'hF3;
            GRN=8'hB0;
            BLU=8'h95;
        end
        1050:
        begin
            RED=8'hEB;
            GRN=8'hAE;
            BLU=8'h91;
        end
        1051:
        begin
            RED=8'hC6;
            GRN=8'h8A;
            BLU=8'h70;
        end
        1052:
        begin
            RED=8'h1A;
            GRN=8'h17;
            BLU=8'h2A;
        end
        1053:
        begin
            RED=8'h1A;
            GRN=8'h17;
            BLU=8'h2A;
        end
        1054:
        begin
            RED=8'h18;
            GRN=8'h15;
            BLU=8'h26;
        end
        1055:
        begin
            RED=8'h17;
            GRN=8'h15;
            BLU=8'h23;
        end
        1056:
        begin
            RED=8'h16;
            GRN=8'h13;
            BLU=8'h24;
        end
        1057:
        begin
            RED=8'h15;
            GRN=8'h13;
            BLU=8'h20;
        end
        1058:
        begin
            RED=8'h12;
            GRN=8'h11;
            BLU=8'h19;
        end
        1059:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        1060:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h15;
        end
        1061:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        1062:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        1063:
        begin
            RED=8'h08;
            GRN=8'h07;
            BLU=8'h0F;
        end
        1088:
        begin
            RED=8'h0C;
            GRN=8'h0B;
            BLU=8'h11;
        end
        1089:
        begin
            RED=8'h0D;
            GRN=8'h10;
            BLU=8'h19;
        end
        1090:
        begin
            RED=8'h14;
            GRN=8'h12;
            BLU=8'h1F;
        end
        1091:
        begin
            RED=8'h14;
            GRN=8'h11;
            BLU=8'h22;
        end
        1092:
        begin
            RED=8'h16;
            GRN=8'h13;
            BLU=8'h24;
        end
        1093:
        begin
            RED=8'h16;
            GRN=8'h15;
            BLU=8'h27;
        end
        1094:
        begin
            RED=8'h19;
            GRN=8'h18;
            BLU=8'h2A;
        end
        1095:
        begin
            RED=8'h19;
            GRN=8'h15;
            BLU=8'h2C;
        end
        1096:
        begin
            RED=8'h1A;
            GRN=8'h16;
            BLU=8'h2D;
        end
        1097:
        begin
            RED=8'h19;
            GRN=8'h15;
            BLU=8'h2C;
        end
        1098:
        begin
            RED=8'h1B;
            GRN=8'h18;
            BLU=8'h2D;
        end
        1099:
        begin
            RED=8'h1C;
            GRN=8'h18;
            BLU=8'h2F;
        end
        1100:
        begin
            RED=8'hE9;
            GRN=8'hB7;
            BLU=8'h9C;
        end
        1101:
        begin
            RED=8'hAB;
            GRN=8'h7E;
            BLU=8'h6B;
        end
        1102:
        begin
            RED=8'hB4;
            GRN=8'h7B;
            BLU=8'h60;
        end
        1103:
        begin
            RED=8'hE8;
            GRN=8'hA6;
            BLU=8'h8C;
        end
        1104:
        begin
            RED=8'hFA;
            GRN=8'hB7;
            BLU=8'h9D;
        end
        1105:
        begin
            RED=8'hFD;
            GRN=8'hB5;
            BLU=8'h9C;
        end
        1106:
        begin
            RED=8'hFF;
            GRN=8'hB5;
            BLU=8'h9C;
        end
        1107:
        begin
            RED=8'hEB;
            GRN=8'hA1;
            BLU=8'h88;
        end
        1108:
        begin
            RED=8'hC5;
            GRN=8'h83;
            BLU=8'h6B;
        end
        1109:
        begin
            RED=8'hF1;
            GRN=8'hA7;
            BLU=8'h8E;
        end
        1110:
        begin
            RED=8'hDC;
            GRN=8'h98;
            BLU=8'h81;
        end
        1111:
        begin
            RED=8'hD9;
            GRN=8'h8D;
            BLU=8'h73;
        end
        1112:
        begin
            RED=8'hEE;
            GRN=8'hA3;
            BLU=8'h8C;
        end
        1113:
        begin
            RED=8'hE8;
            GRN=8'h9C;
            BLU=8'h84;
        end
        1114:
        begin
            RED=8'hDE;
            GRN=8'h9C;
            BLU=8'h86;
        end
        1115:
        begin
            RED=8'hB3;
            GRN=8'h7D;
            BLU=8'h63;
        end
        1116:
        begin
            RED=8'h1C;
            GRN=8'h1B;
            BLU=8'h2D;
        end
        1117:
        begin
            RED=8'h1A;
            GRN=8'h17;
            BLU=8'h2A;
        end
        1118:
        begin
            RED=8'h19;
            GRN=8'h16;
            BLU=8'h29;
        end
        1119:
        begin
            RED=8'h18;
            GRN=8'h15;
            BLU=8'h28;
        end
        1120:
        begin
            RED=8'h17;
            GRN=8'h15;
            BLU=8'h23;
        end
        1121:
        begin
            RED=8'h16;
            GRN=8'h14;
            BLU=8'h21;
        end
        1122:
        begin
            RED=8'h14;
            GRN=8'h13;
            BLU=8'h1B;
        end
        1123:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h1A;
        end
        1124:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h15;
        end
        1125:
        begin
            RED=8'h0C;
            GRN=8'h0B;
            BLU=8'h13;
        end
        1126:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        1127:
        begin
            RED=8'h08;
            GRN=8'h07;
            BLU=8'h0F;
        end
        1152:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h13;
        end
        1153:
        begin
            RED=8'h0F;
            GRN=8'h0D;
            BLU=8'h1A;
        end
        1154:
        begin
            RED=8'h14;
            GRN=8'h12;
            BLU=8'h20;
        end
        1155:
        begin
            RED=8'h15;
            GRN=8'h12;
            BLU=8'h23;
        end
        1156:
        begin
            RED=8'h18;
            GRN=8'h15;
            BLU=8'h28;
        end
        1157:
        begin
            RED=8'h17;
            GRN=8'h16;
            BLU=8'h28;
        end
        1158:
        begin
            RED=8'h1A;
            GRN=8'h17;
            BLU=8'h2C;
        end
        1159:
        begin
            RED=8'h19;
            GRN=8'h15;
            BLU=8'h2C;
        end
        1160:
        begin
            RED=8'h1B;
            GRN=8'h17;
            BLU=8'h2E;
        end
        1161:
        begin
            RED=8'h1B;
            GRN=8'h17;
            BLU=8'h2E;
        end
        1162:
        begin
            RED=8'h1E;
            GRN=8'h1A;
            BLU=8'h33;
        end
        1163:
        begin
            RED=8'h1E;
            GRN=8'h1A;
            BLU=8'h33;
        end
        1164:
        begin
            RED=8'hA6;
            GRN=8'h73;
            BLU=8'h62;
        end
        1165:
        begin
            RED=8'hB7;
            GRN=8'h88;
            BLU=8'h6A;
        end
        1166:
        begin
            RED=8'hAE;
            GRN=8'h7E;
            BLU=8'h68;
        end
        1167:
        begin
            RED=8'hDB;
            GRN=8'h97;
            BLU=8'h80;
        end
        1168:
        begin
            RED=8'hF9;
            GRN=8'hBC;
            BLU=8'hA9;
        end
        1169:
        begin
            RED=8'hF6;
            GRN=8'hA8;
            BLU=8'h91;
        end
        1170:
        begin
            RED=8'hE0;
            GRN=8'h90;
            BLU=8'h77;
        end
        1171:
        begin
            RED=8'hB8;
            GRN=8'h71;
            BLU=8'h5D;
        end
        1172:
        begin
            RED=8'hD1;
            GRN=8'h8F;
            BLU=8'h77;
        end
        1173:
        begin
            RED=8'hEB;
            GRN=8'hA3;
            BLU=8'h8B;
        end
        1174:
        begin
            RED=8'hE0;
            GRN=8'h9E;
            BLU=8'h86;
        end
        1175:
        begin
            RED=8'hD0;
            GRN=8'h85;
            BLU=8'h70;
        end
        1176:
        begin
            RED=8'hAC;
            GRN=8'h5E;
            BLU=8'h47;
        end
        1177:
        begin
            RED=8'hE3;
            GRN=8'h93;
            BLU=8'h7A;
        end
        1178:
        begin
            RED=8'hD2;
            GRN=8'h90;
            BLU=8'h7A;
        end
        1179:
        begin
            RED=8'hA7;
            GRN=8'h7A;
            BLU=8'h65;
        end
        1180:
        begin
            RED=8'h1B;
            GRN=8'h1A;
            BLU=8'h2C;
        end
        1181:
        begin
            RED=8'h1A;
            GRN=8'h19;
            BLU=8'h2B;
        end
        1182:
        begin
            RED=8'h19;
            GRN=8'h18;
            BLU=8'h2A;
        end
        1183:
        begin
            RED=8'h19;
            GRN=8'h16;
            BLU=8'h29;
        end
        1184:
        begin
            RED=8'h16;
            GRN=8'h13;
            BLU=8'h24;
        end
        1185:
        begin
            RED=8'h17;
            GRN=8'h15;
            BLU=8'h23;
        end
        1186:
        begin
            RED=8'h15;
            GRN=8'h13;
            BLU=8'h1E;
        end
        1187:
        begin
            RED=8'h15;
            GRN=8'h13;
            BLU=8'h1E;
        end
        1188:
        begin
            RED=8'h11;
            GRN=8'h0F;
            BLU=8'h1A;
        end
        1189:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h14;
        end
        1190:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        1191:
        begin
            RED=8'h09;
            GRN=8'h08;
            BLU=8'h10;
        end
        1216:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        1217:
        begin
            RED=8'h11;
            GRN=8'h0F;
            BLU=8'h1C;
        end
        1218:
        begin
            RED=8'h14;
            GRN=8'h11;
            BLU=8'h22;
        end
        1219:
        begin
            RED=8'h16;
            GRN=8'h13;
            BLU=8'h26;
        end
        1220:
        begin
            RED=8'h16;
            GRN=8'h14;
            BLU=8'h29;
        end
        1221:
        begin
            RED=8'h17;
            GRN=8'h13;
            BLU=8'h2C;
        end
        1222:
        begin
            RED=8'h1B;
            GRN=8'h17;
            BLU=8'h2E;
        end
        1223:
        begin
            RED=8'h1B;
            GRN=8'h17;
            BLU=8'h30;
        end
        1224:
        begin
            RED=8'h1C;
            GRN=8'h17;
            BLU=8'h35;
        end
        1225:
        begin
            RED=8'h1B;
            GRN=8'h16;
            BLU=8'h34;
        end
        1226:
        begin
            RED=8'h1D;
            GRN=8'h18;
            BLU=8'h36;
        end
        1227:
        begin
            RED=8'h1D;
            GRN=8'h18;
            BLU=8'h36;
        end
        1228:
        begin
            RED=8'h17;
            GRN=8'h0F;
            BLU=8'h26;
        end
        1229:
        begin
            RED=8'hD0;
            GRN=8'h8E;
            BLU=8'h76;
        end
        1230:
        begin
            RED=8'hA1;
            GRN=8'h71;
            BLU=8'h5A;
        end
        1231:
        begin
            RED=8'hBC;
            GRN=8'h7A;
            BLU=8'h62;
        end
        1232:
        begin
            RED=8'hC5;
            GRN=8'h7F;
            BLU=8'h66;
        end
        1233:
        begin
            RED=8'hCD;
            GRN=8'h80;
            BLU=8'h66;
        end
        1234:
        begin
            RED=8'hD0;
            GRN=8'h8E;
            BLU=8'h74;
        end
        1235:
        begin
            RED=8'hD8;
            GRN=8'h9B;
            BLU=8'h89;
        end
        1236:
        begin
            RED=8'hB1;
            GRN=8'h84;
            BLU=8'h71;
        end
        1237:
        begin
            RED=8'h6E;
            GRN=8'h40;
            BLU=8'h33;
        end
        1238:
        begin
            RED=8'h9E;
            GRN=8'h6F;
            BLU=8'h5F;
        end
        1239:
        begin
            RED=8'hC7;
            GRN=8'h92;
            BLU=8'h80;
        end
        1240:
        begin
            RED=8'h9B;
            GRN=8'h6E;
            BLU=8'h59;
        end
        1241:
        begin
            RED=8'hAE;
            GRN=8'h6A;
            BLU=8'h53;
        end
        1242:
        begin
            RED=8'h96;
            GRN=8'h5C;
            BLU=8'h46;
        end
        1243:
        begin
            RED=8'h99;
            GRN=8'h73;
            BLU=8'h60;
        end
        1244:
        begin
            RED=8'h1C;
            GRN=8'h18;
            BLU=8'h2F;
        end
        1245:
        begin
            RED=8'h1A;
            GRN=8'h16;
            BLU=8'h2D;
        end
        1246:
        begin
            RED=8'h1A;
            GRN=8'h17;
            BLU=8'h2C;
        end
        1247:
        begin
            RED=8'h18;
            GRN=8'h16;
            BLU=8'h2B;
        end
        1248:
        begin
            RED=8'h1A;
            GRN=8'h17;
            BLU=8'h2A;
        end
        1249:
        begin
            RED=8'h16;
            GRN=8'h13;
            BLU=8'h24;
        end
        1250:
        begin
            RED=8'h16;
            GRN=8'h14;
            BLU=8'h22;
        end
        1251:
        begin
            RED=8'h15;
            GRN=8'h13;
            BLU=8'h20;
        end
        1252:
        begin
            RED=8'h12;
            GRN=8'h10;
            BLU=8'h1B;
        end
        1253:
        begin
            RED=8'h0F;
            GRN=8'h0E;
            BLU=8'h14;
        end
        1254:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        1255:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        1280:
        begin
            RED=8'h0F;
            GRN=8'h0D;
            BLU=8'h18;
        end
        1281:
        begin
            RED=8'h12;
            GRN=8'h0F;
            BLU=8'h20;
        end
        1282:
        begin
            RED=8'h15;
            GRN=8'h12;
            BLU=8'h23;
        end
        1283:
        begin
            RED=8'h16;
            GRN=8'h13;
            BLU=8'h26;
        end
        1284:
        begin
            RED=8'h16;
            GRN=8'h12;
            BLU=8'h29;
        end
        1285:
        begin
            RED=8'h19;
            GRN=8'h16;
            BLU=8'h2B;
        end
        1286:
        begin
            RED=8'h1A;
            GRN=8'h17;
            BLU=8'h32;
        end
        1287:
        begin
            RED=8'h19;
            GRN=8'h19;
            BLU=8'h33;
        end
        1288:
        begin
            RED=8'h1C;
            GRN=8'h17;
            BLU=8'h37;
        end
        1289:
        begin
            RED=8'h18;
            GRN=8'h15;
            BLU=8'h34;
        end
        1290:
        begin
            RED=8'h1E;
            GRN=8'h1B;
            BLU=8'h3A;
        end
        1291:
        begin
            RED=8'h1C;
            GRN=8'h19;
            BLU=8'h38;
        end
        1292:
        begin
            RED=8'h1B;
            GRN=8'h1A;
            BLU=8'h3A;
        end
        1293:
        begin
            RED=8'h4B;
            GRN=8'h2D;
            BLU=8'h2D;
        end
        1294:
        begin
            RED=8'hAC;
            GRN=8'h79;
            BLU=8'h5C;
        end
        1295:
        begin
            RED=8'hAA;
            GRN=8'h72;
            BLU=8'h59;
        end
        1296:
        begin
            RED=8'hBC;
            GRN=8'h7D;
            BLU=8'h5A;
        end
        1297:
        begin
            RED=8'hC1;
            GRN=8'h8C;
            BLU=8'h6A;
        end
        1298:
        begin
            RED=8'hC5;
            GRN=8'h97;
            BLU=8'h87;
        end
        1299:
        begin
            RED=8'hD2;
            GRN=8'hA5;
            BLU=8'h92;
        end
        1300:
        begin
            RED=8'hC4;
            GRN=8'h8B;
            BLU=8'h7A;
        end
        1301:
        begin
            RED=8'hC1;
            GRN=8'h93;
            BLU=8'h83;
        end
        1302:
        begin
            RED=8'hD1;
            GRN=8'h96;
            BLU=8'h84;
        end
        1303:
        begin
            RED=8'hB5;
            GRN=8'h8D;
            BLU=8'h74;
        end
        1304:
        begin
            RED=8'hAB;
            GRN=8'h79;
            BLU=8'h60;
        end
        1305:
        begin
            RED=8'hC5;
            GRN=8'h7E;
            BLU=8'h60;
        end
        1306:
        begin
            RED=8'hAF;
            GRN=8'h77;
            BLU=8'h60;
        end
        1307:
        begin
            RED=8'h5B;
            GRN=8'h4D;
            BLU=8'h4A;
        end
        1308:
        begin
            RED=8'h1A;
            GRN=8'h18;
            BLU=8'h30;
        end
        1309:
        begin
            RED=8'h1B;
            GRN=8'h18;
            BLU=8'h2D;
        end
        1310:
        begin
            RED=8'h1A;
            GRN=8'h16;
            BLU=8'h2D;
        end
        1311:
        begin
            RED=8'h19;
            GRN=8'h15;
            BLU=8'h2C;
        end
        1312:
        begin
            RED=8'h19;
            GRN=8'h17;
            BLU=8'h2C;
        end
        1313:
        begin
            RED=8'h17;
            GRN=8'h14;
            BLU=8'h27;
        end
        1314:
        begin
            RED=8'h15;
            GRN=8'h12;
            BLU=8'h23;
        end
        1315:
        begin
            RED=8'h14;
            GRN=8'h12;
            BLU=8'h1F;
        end
        1316:
        begin
            RED=8'h11;
            GRN=8'h0F;
            BLU=8'h1A;
        end
        1317:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h17;
        end
        1318:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        1319:
        begin
            RED=8'h09;
            GRN=8'h08;
            BLU=8'h0E;
        end
        1344:
        begin
            RED=8'h11;
            GRN=8'h0F;
            BLU=8'h1C;
        end
        1345:
        begin
            RED=8'h13;
            GRN=8'h10;
            BLU=8'h21;
        end
        1346:
        begin
            RED=8'h14;
            GRN=8'h13;
            BLU=8'h25;
        end
        1347:
        begin
            RED=8'h16;
            GRN=8'h14;
            BLU=8'h29;
        end
        1348:
        begin
            RED=8'h16;
            GRN=8'h13;
            BLU=8'h28;
        end
        1349:
        begin
            RED=8'h1A;
            GRN=8'h16;
            BLU=8'h2F;
        end
        1350:
        begin
            RED=8'h1A;
            GRN=8'h15;
            BLU=8'h33;
        end
        1351:
        begin
            RED=8'h1D;
            GRN=8'h18;
            BLU=8'h36;
        end
        1352:
        begin
            RED=8'h1B;
            GRN=8'h18;
            BLU=8'h37;
        end
        1353:
        begin
            RED=8'h1A;
            GRN=8'h16;
            BLU=8'h39;
        end
        1354:
        begin
            RED=8'h1B;
            GRN=8'h17;
            BLU=8'h3A;
        end
        1355:
        begin
            RED=8'h1A;
            GRN=8'h19;
            BLU=8'h3B;
        end
        1356:
        begin
            RED=8'h1C;
            GRN=8'h18;
            BLU=8'h3B;
        end
        1357:
        begin
            RED=8'h1A;
            GRN=8'h1B;
            BLU=8'h3A;
        end
        1358:
        begin
            RED=8'h96;
            GRN=8'h69;
            BLU=8'h54;
        end
        1359:
        begin
            RED=8'hB2;
            GRN=8'h80;
            BLU=8'h65;
        end
        1360:
        begin
            RED=8'hCA;
            GRN=8'h88;
            BLU=8'h66;
        end
        1361:
        begin
            RED=8'hDD;
            GRN=8'h9C;
            BLU=8'h7C;
        end
        1362:
        begin
            RED=8'hC2;
            GRN=8'h81;
            BLU=8'h6D;
        end
        1363:
        begin
            RED=8'h4D;
            GRN=8'h2D;
            BLU=8'h20;
        end
        1364:
        begin
            RED=8'h8B;
            GRN=8'h5B;
            BLU=8'h44;
        end
        1365:
        begin
            RED=8'h84;
            GRN=8'h46;
            BLU=8'h2D;
        end
        1366:
        begin
            RED=8'hBB;
            GRN=8'hAA;
            BLU=8'h8E;
        end
        1367:
        begin
            RED=8'h9A;
            GRN=8'h4D;
            BLU=8'h45;
        end
        1368:
        begin
            RED=8'hBB;
            GRN=8'h80;
            BLU=8'h62;
        end
        1369:
        begin
            RED=8'hD5;
            GRN=8'h90;
            BLU=8'h71;
        end
        1370:
        begin
            RED=8'hB1;
            GRN=8'h7F;
            BLU=8'h66;
        end
        1371:
        begin
            RED=8'h1E;
            GRN=8'h1A;
            BLU=8'h3B;
        end
        1372:
        begin
            RED=8'h1D;
            GRN=8'h19;
            BLU=8'h34;
        end
        1373:
        begin
            RED=8'h1C;
            GRN=8'h18;
            BLU=8'h33;
        end
        1374:
        begin
            RED=8'h1B;
            GRN=8'h17;
            BLU=8'h2E;
        end
        1375:
        begin
            RED=8'h1A;
            GRN=8'h16;
            BLU=8'h2D;
        end
        1376:
        begin
            RED=8'h1A;
            GRN=8'h17;
            BLU=8'h2C;
        end
        1377:
        begin
            RED=8'h17;
            GRN=8'h16;
            BLU=8'h26;
        end
        1378:
        begin
            RED=8'h16;
            GRN=8'h13;
            BLU=8'h24;
        end
        1379:
        begin
            RED=8'h14;
            GRN=8'h11;
            BLU=8'h22;
        end
        1380:
        begin
            RED=8'h13;
            GRN=8'h11;
            BLU=8'h1E;
        end
        1381:
        begin
            RED=8'h10;
            GRN=8'h0E;
            BLU=8'h1B;
        end
        1382:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        1383:
        begin
            RED=8'h0A;
            GRN=8'h09;
            BLU=8'h11;
        end
        1408:
        begin
            RED=8'h12;
            GRN=8'h10;
            BLU=8'h1D;
        end
        1409:
        begin
            RED=8'h13;
            GRN=8'h10;
            BLU=8'h21;
        end
        1410:
        begin
            RED=8'h14;
            GRN=8'h13;
            BLU=8'h25;
        end
        1411:
        begin
            RED=8'h18;
            GRN=8'h14;
            BLU=8'h2B;
        end
        1412:
        begin
            RED=8'h16;
            GRN=8'h17;
            BLU=8'h2C;
        end
        1413:
        begin
            RED=8'h1A;
            GRN=8'h15;
            BLU=8'h33;
        end
        1414:
        begin
            RED=8'h1A;
            GRN=8'h17;
            BLU=8'h36;
        end
        1415:
        begin
            RED=8'h1C;
            GRN=8'h1B;
            BLU=8'h3A;
        end
        1416:
        begin
            RED=8'h1B;
            GRN=8'h17;
            BLU=8'h38;
        end
        1417:
        begin
            RED=8'h1B;
            GRN=8'h17;
            BLU=8'h3C;
        end
        1418:
        begin
            RED=8'h19;
            GRN=8'h17;
            BLU=8'h3C;
        end
        1419:
        begin
            RED=8'h1C;
            GRN=8'h1A;
            BLU=8'h41;
        end
        1420:
        begin
            RED=8'h1B;
            GRN=8'h1A;
            BLU=8'h39;
        end
        1421:
        begin
            RED=8'h1F;
            GRN=8'h21;
            BLU=8'h20;
        end
        1422:
        begin
            RED=8'h7D;
            GRN=8'h53;
            BLU=8'h3D;
        end
        1423:
        begin
            RED=8'hA5;
            GRN=8'h77;
            BLU=8'h5F;
        end
        1424:
        begin
            RED=8'hB7;
            GRN=8'h7E;
            BLU=8'h60;
        end
        1425:
        begin
            RED=8'hD0;
            GRN=8'h94;
            BLU=8'h70;
        end
        1426:
        begin
            RED=8'hE8;
            GRN=8'hA7;
            BLU=8'h8B;
        end
        1427:
        begin
            RED=8'hD2;
            GRN=8'h8A;
            BLU=8'h71;
        end
        1428:
        begin
            RED=8'hEE;
            GRN=8'h9D;
            BLU=8'h8A;
        end
        1429:
        begin
            RED=8'hE9;
            GRN=8'hAA;
            BLU=8'h9B;
        end
        1430:
        begin
            RED=8'hDA;
            GRN=8'h93;
            BLU=8'h81;
        end
        1431:
        begin
            RED=8'hC6;
            GRN=8'h8C;
            BLU=8'h78;
        end
        1432:
        begin
            RED=8'hDA;
            GRN=8'h9B;
            BLU=8'h7C;
        end
        1433:
        begin
            RED=8'hBF;
            GRN=8'h86;
            BLU=8'h6B;
        end
        1434:
        begin
            RED=8'h93;
            GRN=8'h6F;
            BLU=8'h55;
        end
        1435:
        begin
            RED=8'h1F;
            GRN=8'h1A;
            BLU=8'h38;
        end
        1436:
        begin
            RED=8'h1C;
            GRN=8'h1B;
            BLU=8'h3A;
        end
        1437:
        begin
            RED=8'h1C;
            GRN=8'h17;
            BLU=8'h35;
        end
        1438:
        begin
            RED=8'h1B;
            GRN=8'h16;
            BLU=8'h34;
        end
        1439:
        begin
            RED=8'h1B;
            GRN=8'h17;
            BLU=8'h30;
        end
        1440:
        begin
            RED=8'h1A;
            GRN=8'h17;
            BLU=8'h2A;
        end
        1441:
        begin
            RED=8'h17;
            GRN=8'h13;
            BLU=8'h2A;
        end
        1442:
        begin
            RED=8'h19;
            GRN=8'h16;
            BLU=8'h29;
        end
        1443:
        begin
            RED=8'h16;
            GRN=8'h13;
            BLU=8'h26;
        end
        1444:
        begin
            RED=8'h13;
            GRN=8'h11;
            BLU=8'h1E;
        end
        1445:
        begin
            RED=8'h10;
            GRN=8'h0E;
            BLU=8'h1B;
        end
        1446:
        begin
            RED=8'h0E;
            GRN=8'h0D;
            BLU=8'h15;
        end
        1447:
        begin
            RED=8'h0C;
            GRN=8'h0B;
            BLU=8'h13;
        end
        1472:
        begin
            RED=8'h11;
            GRN=8'h0E;
            BLU=8'h1F;
        end
        1473:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h24;
        end
        1474:
        begin
            RED=8'h15;
            GRN=8'h13;
            BLU=8'h29;
        end
        1475:
        begin
            RED=8'h18;
            GRN=8'h14;
            BLU=8'h2B;
        end
        1476:
        begin
            RED=8'h19;
            GRN=8'h15;
            BLU=8'h30;
        end
        1477:
        begin
            RED=8'h19;
            GRN=8'h14;
            BLU=8'h34;
        end
        1478:
        begin
            RED=8'h19;
            GRN=8'h18;
            BLU=8'h38;
        end
        1479:
        begin
            RED=8'h1B;
            GRN=8'h17;
            BLU=8'h3C;
        end
        1480:
        begin
            RED=8'h19;
            GRN=8'h17;
            BLU=8'h3C;
        end
        1481:
        begin
            RED=8'h1A;
            GRN=8'h18;
            BLU=8'h3F;
        end
        1482:
        begin
            RED=8'h1B;
            GRN=8'h19;
            BLU=8'h40;
        end
        1483:
        begin
            RED=8'h1C;
            GRN=8'h1A;
            BLU=8'h41;
        end
        1484:
        begin
            RED=8'h1B;
            GRN=8'h1B;
            BLU=8'h37;
        end
        1485:
        begin
            RED=8'h12;
            GRN=8'h13;
            BLU=8'h0B;
        end
        1486:
        begin
            RED=8'hE4;
            GRN=8'hE3;
            BLU=8'hDF;
        end
        1487:
        begin
            RED=8'h74;
            GRN=8'h4F;
            BLU=8'h3D;
        end
        1488:
        begin
            RED=8'hA9;
            GRN=8'h7A;
            BLU=8'h5E;
        end
        1489:
        begin
            RED=8'hD5;
            GRN=8'h94;
            BLU=8'h76;
        end
        1490:
        begin
            RED=8'hEE;
            GRN=8'hAE;
            BLU=8'h92;
        end
        1491:
        begin
            RED=8'hD3;
            GRN=8'h95;
            BLU=8'h7E;
        end
        1492:
        begin
            RED=8'hC6;
            GRN=8'h88;
            BLU=8'h71;
        end
        1493:
        begin
            RED=8'hDA;
            GRN=8'h98;
            BLU=8'h82;
        end
        1494:
        begin
            RED=8'hC9;
            GRN=8'h8B;
            BLU=8'h74;
        end
        1495:
        begin
            RED=8'hD7;
            GRN=8'h9B;
            BLU=8'h81;
        end
        1496:
        begin
            RED=8'hD9;
            GRN=8'h9E;
            BLU=8'h80;
        end
        1497:
        begin
            RED=8'h95;
            GRN=8'h67;
            BLU=8'h50;
        end
        1498:
        begin
            RED=8'h1D;
            GRN=8'h1E;
            BLU=8'h3C;
        end
        1499:
        begin
            RED=8'h1F;
            GRN=8'h19;
            BLU=8'h3F;
        end
        1500:
        begin
            RED=8'h1C;
            GRN=8'h19;
            BLU=8'h38;
        end
        1501:
        begin
            RED=8'h1B;
            GRN=8'h18;
            BLU=8'h37;
        end
        1502:
        begin
            RED=8'h1C;
            GRN=8'h17;
            BLU=8'h35;
        end
        1503:
        begin
            RED=8'h1A;
            GRN=8'h16;
            BLU=8'h2F;
        end
        1504:
        begin
            RED=8'h1A;
            GRN=8'h16;
            BLU=8'h2F;
        end
        1505:
        begin
            RED=8'h17;
            GRN=8'h13;
            BLU=8'h2A;
        end
        1506:
        begin
            RED=8'h17;
            GRN=8'h15;
            BLU=8'h2A;
        end
        1507:
        begin
            RED=8'h16;
            GRN=8'h13;
            BLU=8'h26;
        end
        1508:
        begin
            RED=8'h13;
            GRN=8'h11;
            BLU=8'h1F;
        end
        1509:
        begin
            RED=8'h11;
            GRN=8'h0F;
            BLU=8'h1C;
        end
        1510:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        1511:
        begin
            RED=8'h0B;
            GRN=8'h0A;
            BLU=8'h12;
        end
        1536:
        begin
            RED=8'h11;
            GRN=8'h0F;
            BLU=8'h1D;
        end
        1537:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h24;
        end
        1538:
        begin
            RED=8'h16;
            GRN=8'h12;
            BLU=8'h29;
        end
        1539:
        begin
            RED=8'h17;
            GRN=8'h14;
            BLU=8'h2F;
        end
        1540:
        begin
            RED=8'h16;
            GRN=8'h15;
            BLU=8'h34;
        end
        1541:
        begin
            RED=8'h17;
            GRN=8'h16;
            BLU=8'h35;
        end
        1542:
        begin
            RED=8'h19;
            GRN=8'h17;
            BLU=8'h3C;
        end
        1543:
        begin
            RED=8'h18;
            GRN=8'h17;
            BLU=8'h39;
        end
        1544:
        begin
            RED=8'h19;
            GRN=8'h17;
            BLU=8'h3E;
        end
        1545:
        begin
            RED=8'h19;
            GRN=8'h17;
            BLU=8'h3F;
        end
        1546:
        begin
            RED=8'h1A;
            GRN=8'h17;
            BLU=8'h42;
        end
        1547:
        begin
            RED=8'h1A;
            GRN=8'h18;
            BLU=8'h40;
        end
        1548:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h23;
        end
        1549:
        begin
            RED=8'h1B;
            GRN=8'h19;
            BLU=8'h1A;
        end
        1550:
        begin
            RED=8'hDA;
            GRN=8'hD9;
            BLU=8'hE1;
        end
        1551:
        begin
            RED=8'hA2;
            GRN=8'h75;
            BLU=8'h5E;
        end
        1552:
        begin
            RED=8'h73;
            GRN=8'h49;
            BLU=8'h3D;
        end
        1553:
        begin
            RED=8'hAC;
            GRN=8'h76;
            BLU=8'h5A;
        end
        1554:
        begin
            RED=8'hC7;
            GRN=8'h8F;
            BLU=8'h76;
        end
        1555:
        begin
            RED=8'hF6;
            GRN=8'hB7;
            BLU=8'h98;
        end
        1556:
        begin
            RED=8'hE9;
            GRN=8'hA6;
            BLU=8'h8C;
        end
        1557:
        begin
            RED=8'hF1;
            GRN=8'hAA;
            BLU=8'h94;
        end
        1558:
        begin
            RED=8'hEC;
            GRN=8'hA2;
            BLU=8'h89;
        end
        1559:
        begin
            RED=8'hE5;
            GRN=8'h9D;
            BLU=8'h84;
        end
        1560:
        begin
            RED=8'hAD;
            GRN=8'h7E;
            BLU=8'h62;
        end
        1561:
        begin
            RED=8'h23;
            GRN=8'h20;
            BLU=8'h1B;
        end
        1562:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h25;
        end
        1563:
        begin
            RED=8'h25;
            GRN=8'h25;
            BLU=8'h27;
        end
        1564:
        begin
            RED=8'h26;
            GRN=8'h26;
            BLU=8'h26;
        end
        1565:
        begin
            RED=8'h25;
            GRN=8'h25;
            BLU=8'h25;
        end
        1566:
        begin
            RED=8'h27;
            GRN=8'h27;
            BLU=8'h27;
        end
        1567:
        begin
            RED=8'h24;
            GRN=8'h24;
            BLU=8'h26;
        end
        1568:
        begin
            RED=8'h1A;
            GRN=8'h16;
            BLU=8'h2F;
        end
        1569:
        begin
            RED=8'h19;
            GRN=8'h16;
            BLU=8'h2B;
        end
        1570:
        begin
            RED=8'h17;
            GRN=8'h15;
            BLU=8'h2A;
        end
        1571:
        begin
            RED=8'h14;
            GRN=8'h12;
            BLU=8'h27;
        end
        1572:
        begin
            RED=8'h12;
            GRN=8'h10;
            BLU=8'h1D;
        end
        1573:
        begin
            RED=8'h12;
            GRN=8'h10;
            BLU=8'h1D;
        end
        1574:
        begin
            RED=8'h10;
            GRN=8'h0E;
            BLU=8'h1B;
        end
        1575:
        begin
            RED=8'h0C;
            GRN=8'h0B;
            BLU=8'h13;
        end
        1600:
        begin
            RED=8'h10;
            GRN=8'h0F;
            BLU=8'h1F;
        end
        1601:
        begin
            RED=8'h14;
            GRN=8'h11;
            BLU=8'h26;
        end
        1602:
        begin
            RED=8'h17;
            GRN=8'h13;
            BLU=8'h2C;
        end
        1603:
        begin
            RED=8'h16;
            GRN=8'h13;
            BLU=8'h30;
        end
        1604:
        begin
            RED=8'h17;
            GRN=8'h16;
            BLU=8'h35;
        end
        1605:
        begin
            RED=8'h1A;
            GRN=8'h16;
            BLU=8'h39;
        end
        1606:
        begin
            RED=8'h19;
            GRN=8'h17;
            BLU=8'h3E;
        end
        1607:
        begin
            RED=8'h15;
            GRN=8'h17;
            BLU=8'h3E;
        end
        1608:
        begin
            RED=8'h18;
            GRN=8'h16;
            BLU=8'h3B;
        end
        1609:
        begin
            RED=8'h18;
            GRN=8'h16;
            BLU=8'h3D;
        end
        1610:
        begin
            RED=8'h21;
            GRN=8'h1D;
            BLU=8'h38;
        end
        1611:
        begin
            RED=8'h25;
            GRN=8'h25;
            BLU=8'h27;
        end
        1612:
        begin
            RED=8'h26;
            GRN=8'h26;
            BLU=8'h26;
        end
        1613:
        begin
            RED=8'h24;
            GRN=8'h24;
            BLU=8'h24;
        end
        1614:
        begin
            RED=8'hF0;
            GRN=8'hF5;
            BLU=8'hF8;
        end
        1615:
        begin
            RED=8'hDE;
            GRN=8'hE3;
            BLU=8'hE7;
        end
        1616:
        begin
            RED=8'h8F;
            GRN=8'h64;
            BLU=8'h51;
        end
        1617:
        begin
            RED=8'h68;
            GRN=8'h4B;
            BLU=8'h3D;
        end
        1618:
        begin
            RED=8'h73;
            GRN=8'h50;
            BLU=8'h3D;
        end
        1619:
        begin
            RED=8'hC3;
            GRN=8'h87;
            BLU=8'h6B;
        end
        1620:
        begin
            RED=8'hDA;
            GRN=8'h9A;
            BLU=8'h7F;
        end
        1621:
        begin
            RED=8'hD0;
            GRN=8'h8F;
            BLU=8'h71;
        end
        1622:
        begin
            RED=8'hDB;
            GRN=8'h95;
            BLU=8'h7B;
        end
        1623:
        begin
            RED=8'hC4;
            GRN=8'h8B;
            BLU=8'h6E;
        end
        1624:
        begin
            RED=8'h6E;
            GRN=8'h52;
            BLU=8'h46;
        end
        1625:
        begin
            RED=8'h1E;
            GRN=8'h1E;
            BLU=8'h1C;
        end
        1626:
        begin
            RED=8'h1F;
            GRN=8'h1F;
            BLU=8'h1F;
        end
        1627:
        begin
            RED=8'h22;
            GRN=8'h22;
            BLU=8'h24;
        end
        1628:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h23;
        end
        1629:
        begin
            RED=8'h24;
            GRN=8'h24;
            BLU=8'h24;
        end
        1630:
        begin
            RED=8'h24;
            GRN=8'h24;
            BLU=8'h26;
        end
        1631:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h25;
        end
        1632:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h25;
        end
        1633:
        begin
            RED=8'h1C;
            GRN=8'h1A;
            BLU=8'h25;
        end
        1634:
        begin
            RED=8'h17;
            GRN=8'h13;
            BLU=8'h2A;
        end
        1635:
        begin
            RED=8'h16;
            GRN=8'h14;
            BLU=8'h29;
        end
        1636:
        begin
            RED=8'h15;
            GRN=8'h12;
            BLU=8'h23;
        end
        1637:
        begin
            RED=8'h11;
            GRN=8'h0F;
            BLU=8'h1D;
        end
        1638:
        begin
            RED=8'h10;
            GRN=8'h0E;
            BLU=8'h1B;
        end
        1639:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        1664:
        begin
            RED=8'h13;
            GRN=8'h11;
            BLU=8'h26;
        end
        1665:
        begin
            RED=8'h11;
            GRN=8'h0F;
            BLU=8'h24;
        end
        1666:
        begin
            RED=8'h15;
            GRN=8'h13;
            BLU=8'h2B;
        end
        1667:
        begin
            RED=8'h17;
            GRN=8'h14;
            BLU=8'h33;
        end
        1668:
        begin
            RED=8'h19;
            GRN=8'h15;
            BLU=8'h38;
        end
        1669:
        begin
            RED=8'h17;
            GRN=8'h15;
            BLU=8'h3A;
        end
        1670:
        begin
            RED=8'h18;
            GRN=8'h16;
            BLU=8'h3D;
        end
        1671:
        begin
            RED=8'h18;
            GRN=8'h16;
            BLU=8'h3D;
        end
        1672:
        begin
            RED=8'h19;
            GRN=8'h16;
            BLU=8'h41;
        end
        1673:
        begin
            RED=8'h25;
            GRN=8'h26;
            BLU=8'h28;
        end
        1674:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        1675:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h20;
        end
        1676:
        begin
            RED=8'h26;
            GRN=8'h26;
            BLU=8'h26;
        end
        1677:
        begin
            RED=8'h26;
            GRN=8'h26;
            BLU=8'h26;
        end
        1678:
        begin
            RED=8'h1B;
            GRN=8'h1C;
            BLU=8'h1E;
        end
        1679:
        begin
            RED=8'hE9;
            GRN=8'hEC;
            BLU=8'hF1;
        end
        1680:
        begin
            RED=8'hE6;
            GRN=8'hE7;
            BLU=8'hE9;
        end
        1681:
        begin
            RED=8'h80;
            GRN=8'h56;
            BLU=8'h3D;
        end
        1682:
        begin
            RED=8'h6A;
            GRN=8'h4E;
            BLU=8'h42;
        end
        1683:
        begin
            RED=8'h6D;
            GRN=8'h56;
            BLU=8'h4E;
        end
        1684:
        begin
            RED=8'h6B;
            GRN=8'h55;
            BLU=8'h47;
        end
        1685:
        begin
            RED=8'h68;
            GRN=8'h4C;
            BLU=8'h40;
        end
        1686:
        begin
            RED=8'h72;
            GRN=8'h56;
            BLU=8'h48;
        end
        1687:
        begin
            RED=8'h81;
            GRN=8'h68;
            BLU=8'h54;
        end
        1688:
        begin
            RED=8'h5B;
            GRN=8'h3E;
            BLU=8'h30;
        end
        1689:
        begin
            RED=8'h0F;
            GRN=8'h0F;
            BLU=8'h0D;
        end
        1690:
        begin
            RED=8'h1E;
            GRN=8'h1E;
            BLU=8'h1E;
        end
        1691:
        begin
            RED=8'h1F;
            GRN=8'h1F;
            BLU=8'h1F;
        end
        1692:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h25;
        end
        1693:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h25;
        end
        1694:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h25;
        end
        1695:
        begin
            RED=8'h21;
            GRN=8'h21;
            BLU=8'h23;
        end
        1696:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h22;
        end
        1697:
        begin
            RED=8'h21;
            GRN=8'h21;
            BLU=8'h23;
        end
        1698:
        begin
            RED=8'h12;
            GRN=8'h12;
            BLU=8'h10;
        end
        1699:
        begin
            RED=8'h15;
            GRN=8'h13;
            BLU=8'h28;
        end
        1700:
        begin
            RED=8'h14;
            GRN=8'h11;
            BLU=8'h22;
        end
        1701:
        begin
            RED=8'h12;
            GRN=8'h10;
            BLU=8'h1E;
        end
        1702:
        begin
            RED=8'h11;
            GRN=8'h0F;
            BLU=8'h1C;
        end
        1703:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        1728:
        begin
            RED=8'h12;
            GRN=8'h0E;
            BLU=8'h25;
        end
        1729:
        begin
            RED=8'h14;
            GRN=8'h12;
            BLU=8'h2A;
        end
        1730:
        begin
            RED=8'h14;
            GRN=8'h14;
            BLU=8'h30;
        end
        1731:
        begin
            RED=8'h15;
            GRN=8'h14;
            BLU=8'h34;
        end
        1732:
        begin
            RED=8'h17;
            GRN=8'h16;
            BLU=8'h38;
        end
        1733:
        begin
            RED=8'h18;
            GRN=8'h16;
            BLU=8'h3D;
        end
        1734:
        begin
            RED=8'h19;
            GRN=8'h17;
            BLU=8'h3E;
        end
        1735:
        begin
            RED=8'h1A;
            GRN=8'h18;
            BLU=8'h3D;
        end
        1736:
        begin
            RED=8'h27;
            GRN=8'h27;
            BLU=8'h25;
        end
        1737:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h2A;
        end
        1738:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        1739:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h23;
        end
        1740:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        1741:
        begin
            RED=8'h27;
            GRN=8'h27;
            BLU=8'h27;
        end
        1742:
        begin
            RED=8'h27;
            GRN=8'h27;
            BLU=8'h29;
        end
        1743:
        begin
            RED=8'hE9;
            GRN=8'hEA;
            BLU=8'hEF;
        end
        1744:
        begin
            RED=8'hED;
            GRN=8'hF2;
            BLU=8'hF6;
        end
        1745:
        begin
            RED=8'hE9;
            GRN=8'hEB;
            BLU=8'hEA;
        end
        1746:
        begin
            RED=8'h8F;
            GRN=8'h7E;
            BLU=8'h6C;
        end
        1747:
        begin
            RED=8'h78;
            GRN=8'h59;
            BLU=8'h45;
        end
        1748:
        begin
            RED=8'h74;
            GRN=8'h56;
            BLU=8'h3E;
        end
        1749:
        begin
            RED=8'h77;
            GRN=8'h58;
            BLU=8'h44;
        end
        1750:
        begin
            RED=8'h7C;
            GRN=8'h59;
            BLU=8'h45;
        end
        1751:
        begin
            RED=8'h8E;
            GRN=8'h72;
            BLU=8'h5C;
        end
        1752:
        begin
            RED=8'hEC;
            GRN=8'hE6;
            BLU=8'hE6;
        end
        1753:
        begin
            RED=8'h24;
            GRN=8'h24;
            BLU=8'h22;
        end
        1754:
        begin
            RED=8'h1C;
            GRN=8'h1C;
            BLU=8'h1C;
        end
        1755:
        begin
            RED=8'h1F;
            GRN=8'h1F;
            BLU=8'h1F;
        end
        1756:
        begin
            RED=8'h22;
            GRN=8'h22;
            BLU=8'h24;
        end
        1757:
        begin
            RED=8'h21;
            GRN=8'h21;
            BLU=8'h23;
        end
        1758:
        begin
            RED=8'h22;
            GRN=8'h22;
            BLU=8'h24;
        end
        1759:
        begin
            RED=8'h22;
            GRN=8'h22;
            BLU=8'h24;
        end
        1760:
        begin
            RED=8'h21;
            GRN=8'h21;
            BLU=8'h23;
        end
        1761:
        begin
            RED=8'h1E;
            GRN=8'h1E;
            BLU=8'h1E;
        end
        1762:
        begin
            RED=8'h1A;
            GRN=8'h1A;
            BLU=8'h1A;
        end
        1763:
        begin
            RED=8'h1B;
            GRN=8'h1B;
            BLU=8'h1B;
        end
        1764:
        begin
            RED=8'h15;
            GRN=8'h12;
            BLU=8'h27;
        end
        1765:
        begin
            RED=8'h13;
            GRN=8'h11;
            BLU=8'h1F;
        end
        1766:
        begin
            RED=8'h10;
            GRN=8'h0E;
            BLU=8'h1B;
        end
        1767:
        begin
            RED=8'h0E;
            GRN=8'h0C;
            BLU=8'h17;
        end
        1792:
        begin
            RED=8'h12;
            GRN=8'h0E;
            BLU=8'h25;
        end
        1793:
        begin
            RED=8'h11;
            GRN=8'h12;
            BLU=8'h27;
        end
        1794:
        begin
            RED=8'h16;
            GRN=8'h12;
            BLU=8'h33;
        end
        1795:
        begin
            RED=8'h18;
            GRN=8'h15;
            BLU=8'h34;
        end
        1796:
        begin
            RED=8'h18;
            GRN=8'h17;
            BLU=8'h41;
        end
        1797:
        begin
            RED=8'h11;
            GRN=8'h14;
            BLU=8'h35;
        end
        1798:
        begin
            RED=8'h23;
            GRN=8'h24;
            BLU=8'h1F;
        end
        1799:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        1800:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        1801:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        1802:
        begin
            RED=8'h25;
            GRN=8'h25;
            BLU=8'h25;
        end
        1803:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h23;
        end
        1804:
        begin
            RED=8'h2B;
            GRN=8'h2B;
            BLU=8'h2D;
        end
        1805:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2C;
        end
        1806:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        1807:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        1808:
        begin
            RED=8'hE5;
            GRN=8'hE8;
            BLU=8'hED;
        end
        1809:
        begin
            RED=8'hEF;
            GRN=8'hF3;
            BLU=8'hF6;
        end
        1810:
        begin
            RED=8'hF0;
            GRN=8'hF4;
            BLU=8'hF7;
        end
        1811:
        begin
            RED=8'hDB;
            GRN=8'hDB;
            BLU=8'hDD;
        end
        1812:
        begin
            RED=8'hA9;
            GRN=8'h87;
            BLU=8'h6E;
        end
        1813:
        begin
            RED=8'h9D;
            GRN=8'h78;
            BLU=8'h65;
        end
        1814:
        begin
            RED=8'h93;
            GRN=8'h6D;
            BLU=8'h5A;
        end
        1815:
        begin
            RED=8'h9A;
            GRN=8'h70;
            BLU=8'h58;
        end
        1816:
        begin
            RED=8'hF1;
            GRN=8'hF5;
            BLU=8'hF6;
        end
        1817:
        begin
            RED=8'h51;
            GRN=8'h53;
            BLU=8'h4E;
        end
        1818:
        begin
            RED=8'h1D;
            GRN=8'h1D;
            BLU=8'h1D;
        end
        1819:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h20;
        end
        1820:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h22;
        end
        1821:
        begin
            RED=8'h1F;
            GRN=8'h1F;
            BLU=8'h21;
        end
        1822:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h22;
        end
        1823:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h22;
        end
        1824:
        begin
            RED=8'h21;
            GRN=8'h21;
            BLU=8'h23;
        end
        1825:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h20;
        end
        1826:
        begin
            RED=8'h1B;
            GRN=8'h1B;
            BLU=8'h1B;
        end
        1827:
        begin
            RED=8'h19;
            GRN=8'h19;
            BLU=8'h19;
        end
        1828:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h24;
        end
        1829:
        begin
            RED=8'h13;
            GRN=8'h10;
            BLU=8'h21;
        end
        1830:
        begin
            RED=8'h10;
            GRN=8'h0D;
            BLU=8'h1E;
        end
        1831:
        begin
            RED=8'h0F;
            GRN=8'h0D;
            BLU=8'h1A;
        end
        1856:
        begin
            RED=8'h13;
            GRN=8'h10;
            BLU=8'h25;
        end
        1857:
        begin
            RED=8'h12;
            GRN=8'h12;
            BLU=8'h2A;
        end
        1858:
        begin
            RED=8'h14;
            GRN=8'h13;
            BLU=8'h33;
        end
        1859:
        begin
            RED=8'h15;
            GRN=8'h13;
            BLU=8'h38;
        end
        1860:
        begin
            RED=8'h19;
            GRN=8'h12;
            BLU=8'h3C;
        end
        1861:
        begin
            RED=8'h21;
            GRN=8'h21;
            BLU=8'h23;
        end
        1862:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        1863:
        begin
            RED=8'h2B;
            GRN=8'h2B;
            BLU=8'h2D;
        end
        1864:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h29;
        end
        1865:
        begin
            RED=8'h27;
            GRN=8'h27;
            BLU=8'h27;
        end
        1866:
        begin
            RED=8'h27;
            GRN=8'h27;
            BLU=8'h27;
        end
        1867:
        begin
            RED=8'h26;
            GRN=8'h26;
            BLU=8'h26;
        end
        1868:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h23;
        end
        1869:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        1870:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2A;
        end
        1871:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h29;
        end
        1872:
        begin
            RED=8'h1B;
            GRN=8'h1D;
            BLU=8'h1A;
        end
        1873:
        begin
            RED=8'hDD;
            GRN=8'hE2;
            BLU=8'hE5;
        end
        1874:
        begin
            RED=8'hEC;
            GRN=8'hF0;
            BLU=8'hF3;
        end
        1875:
        begin
            RED=8'hF8;
            GRN=8'hFC;
            BLU=8'hFD;
        end
        1876:
        begin
            RED=8'hF4;
            GRN=8'hF4;
            BLU=8'hF6;
        end
        1877:
        begin
            RED=8'hE9;
            GRN=8'hDF;
            BLU=8'hD3;
        end
        1878:
        begin
            RED=8'hA2;
            GRN=8'h78;
            BLU=8'h60;
        end
        1879:
        begin
            RED=8'hFE;
            GRN=8'hFF;
            BLU=8'hFD;
        end
        1880:
        begin
            RED=8'hFA;
            GRN=8'hFF;
            BLU=8'hFB;
        end
        1881:
        begin
            RED=8'h68;
            GRN=8'h67;
            BLU=8'h65;
        end
        1882:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h20;
        end
        1883:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h20;
        end
        1884:
        begin
            RED=8'h21;
            GRN=8'h21;
            BLU=8'h23;
        end
        1885:
        begin
            RED=8'h1F;
            GRN=8'h1F;
            BLU=8'h21;
        end
        1886:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h22;
        end
        1887:
        begin
            RED=8'h21;
            GRN=8'h21;
            BLU=8'h23;
        end
        1888:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h22;
        end
        1889:
        begin
            RED=8'h1F;
            GRN=8'h1F;
            BLU=8'h1F;
        end
        1890:
        begin
            RED=8'h19;
            GRN=8'h19;
            BLU=8'h19;
        end
        1891:
        begin
            RED=8'h18;
            GRN=8'h18;
            BLU=8'h18;
        end
        1892:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h24;
        end
        1893:
        begin
            RED=8'h13;
            GRN=8'h10;
            BLU=8'h21;
        end
        1894:
        begin
            RED=8'h10;
            GRN=8'h0E;
            BLU=8'h1B;
        end
        1895:
        begin
            RED=8'h0E;
            GRN=8'h0C;
            BLU=8'h19;
        end
        1920:
        begin
            RED=8'h13;
            GRN=8'h0F;
            BLU=8'h26;
        end
        1921:
        begin
            RED=8'h14;
            GRN=8'h12;
            BLU=8'h28;
        end
        1922:
        begin
            RED=8'h15;
            GRN=8'h14;
            BLU=8'h34;
        end
        1923:
        begin
            RED=8'h1E;
            GRN=8'h1B;
            BLU=8'h2C;
        end
        1924:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h23;
        end
        1925:
        begin
            RED=8'h25;
            GRN=8'h25;
            BLU=8'h25;
        end
        1926:
        begin
            RED=8'h22;
            GRN=8'h22;
            BLU=8'h22;
        end
        1927:
        begin
            RED=8'h27;
            GRN=8'h27;
            BLU=8'h27;
        end
        1928:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        1929:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2C;
        end
        1930:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        1931:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2C;
        end
        1932:
        begin
            RED=8'h24;
            GRN=8'h24;
            BLU=8'h24;
        end
        1933:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h29;
        end
        1934:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2C;
        end
        1935:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        1936:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2A;
        end
        1937:
        begin
            RED=8'hE4;
            GRN=8'hE6;
            BLU=8'hE5;
        end
        1938:
        begin
            RED=8'hE2;
            GRN=8'hE6;
            BLU=8'hE9;
        end
        1939:
        begin
            RED=8'hED;
            GRN=8'hF1;
            BLU=8'hF4;
        end
        1940:
        begin
            RED=8'hFF;
            GRN=8'hFF;
            BLU=8'hFF;
        end
        1941:
        begin
            RED=8'hFE;
            GRN=8'hFD;
            BLU=8'hFB;
        end
        1942:
        begin
            RED=8'h45;
            GRN=8'h1B;
            BLU=8'h29;
        end
        1943:
        begin
            RED=8'h7A;
            GRN=8'h3B;
            BLU=8'h36;
        end
        1944:
        begin
            RED=8'h82;
            GRN=8'h76;
            BLU=8'h78;
        end
        1945:
        begin
            RED=8'hEA;
            GRN=8'hEC;
            BLU=8'hE7;
        end
        1946:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h23;
        end
        1947:
        begin
            RED=8'h1E;
            GRN=8'h1E;
            BLU=8'h1E;
        end
        1948:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h22;
        end
        1949:
        begin
            RED=8'h21;
            GRN=8'h21;
            BLU=8'h23;
        end
        1950:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h22;
        end
        1951:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h22;
        end
        1952:
        begin
            RED=8'h1F;
            GRN=8'h1F;
            BLU=8'h21;
        end
        1953:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h20;
        end
        1954:
        begin
            RED=8'h1A;
            GRN=8'h1A;
            BLU=8'h1A;
        end
        1955:
        begin
            RED=8'h10;
            GRN=8'h10;
            BLU=8'h10;
        end
        1956:
        begin
            RED=8'h15;
            GRN=8'h16;
            BLU=8'h1B;
        end
        1957:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h24;
        end
        1958:
        begin
            RED=8'h11;
            GRN=8'h0F;
            BLU=8'h1D;
        end
        1959:
        begin
            RED=8'h0D;
            GRN=8'h0B;
            BLU=8'h18;
        end
        1984:
        begin
            RED=8'h12;
            GRN=8'h10;
            BLU=8'h26;
        end
        1985:
        begin
            RED=8'h15;
            GRN=8'h12;
            BLU=8'h2F;
        end
        1986:
        begin
            RED=8'h1C;
            GRN=8'h1C;
            BLU=8'h1E;
        end
        1987:
        begin
            RED=8'h21;
            GRN=8'h21;
            BLU=8'h21;
        end
        1988:
        begin
            RED=8'h24;
            GRN=8'h24;
            BLU=8'h24;
        end
        1989:
        begin
            RED=8'h25;
            GRN=8'h25;
            BLU=8'h25;
        end
        1990:
        begin
            RED=8'h26;
            GRN=8'h26;
            BLU=8'h26;
        end
        1991:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h29;
        end
        1992:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        1993:
        begin
            RED=8'h2B;
            GRN=8'h2B;
            BLU=8'h2D;
        end
        1994:
        begin
            RED=8'h2C;
            GRN=8'h2C;
            BLU=8'h2E;
        end
        1995:
        begin
            RED=8'h2B;
            GRN=8'h2B;
            BLU=8'h2D;
        end
        1996:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        1997:
        begin
            RED=8'h1D;
            GRN=8'h1D;
            BLU=8'h1D;
        end
        1998:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        1999:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        2000:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2A;
        end
        2001:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2002:
        begin
            RED=8'hE1;
            GRN=8'hE1;
            BLU=8'hDF;
        end
        2003:
        begin
            RED=8'hE2;
            GRN=8'hE6;
            BLU=8'hE7;
        end
        2004:
        begin
            RED=8'hF6;
            GRN=8'hF8;
            BLU=8'hF7;
        end
        2005:
        begin
            RED=8'hFF;
            GRN=8'hFE;
            BLU=8'hF9;
        end
        2006:
        begin
            RED=8'hA6;
            GRN=8'h40;
            BLU=8'h31;
        end
        2007:
        begin
            RED=8'hA5;
            GRN=8'h8B;
            BLU=8'hA4;
        end
        2008:
        begin
            RED=8'h4A;
            GRN=8'h38;
            BLU=8'h34;
        end
        2009:
        begin
            RED=8'hDF;
            GRN=8'hE8;
            BLU=8'hE5;
        end
        2010:
        begin
            RED=8'h25;
            GRN=8'h25;
            BLU=8'h25;
        end
        2011:
        begin
            RED=8'h24;
            GRN=8'h24;
            BLU=8'h24;
        end
        2012:
        begin
            RED=8'h1F;
            GRN=8'h1F;
            BLU=8'h21;
        end
        2013:
        begin
            RED=8'h22;
            GRN=8'h22;
            BLU=8'h24;
        end
        2014:
        begin
            RED=8'h21;
            GRN=8'h21;
            BLU=8'h23;
        end
        2015:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h22;
        end
        2016:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h22;
        end
        2017:
        begin
            RED=8'h1F;
            GRN=8'h1F;
            BLU=8'h1F;
        end
        2018:
        begin
            RED=8'h1D;
            GRN=8'h1D;
            BLU=8'h1D;
        end
        2019:
        begin
            RED=8'h0B;
            GRN=8'h0B;
            BLU=8'h0B;
        end
        2020:
        begin
            RED=8'h15;
            GRN=8'h15;
            BLU=8'h17;
        end
        2021:
        begin
            RED=8'h13;
            GRN=8'h12;
            BLU=8'h24;
        end
        2022:
        begin
            RED=8'h10;
            GRN=8'h0D;
            BLU=8'h1E;
        end
        2023:
        begin
            RED=8'h0D;
            GRN=8'h0B;
            BLU=8'h16;
        end
        2048:
        begin
            RED=8'h13;
            GRN=8'h11;
            BLU=8'h27;
        end
        2049:
        begin
            RED=8'h18;
            GRN=8'h18;
            BLU=8'h1A;
        end
        2050:
        begin
            RED=8'h1F;
            GRN=8'h1F;
            BLU=8'h1F;
        end
        2051:
        begin
            RED=8'h21;
            GRN=8'h21;
            BLU=8'h21;
        end
        2052:
        begin
            RED=8'h25;
            GRN=8'h25;
            BLU=8'h25;
        end
        2053:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2054:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2C;
        end
        2055:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2C;
        end
        2056:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2A;
        end
        2057:
        begin
            RED=8'h2B;
            GRN=8'h2B;
            BLU=8'h2D;
        end
        2058:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h2A;
        end
        2059:
        begin
            RED=8'h2B;
            GRN=8'h2B;
            BLU=8'h2D;
        end
        2060:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        2061:
        begin
            RED=8'h27;
            GRN=8'h27;
            BLU=8'h29;
        end
        2062:
        begin
            RED=8'h27;
            GRN=8'h27;
            BLU=8'h27;
        end
        2063:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h29;
        end
        2064:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2065:
        begin
            RED=8'h2B;
            GRN=8'h2B;
            BLU=8'h2B;
        end
        2066:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2A;
        end
        2067:
        begin
            RED=8'hE5;
            GRN=8'hE6;
            BLU=8'hE8;
        end
        2068:
        begin
            RED=8'hF2;
            GRN=8'hF6;
            BLU=8'hF7;
        end
        2069:
        begin
            RED=8'h68;
            GRN=8'h5E;
            BLU=8'h5D;
        end
        2070:
        begin
            RED=8'h4B;
            GRN=8'h23;
            BLU=8'h2C;
        end
        2071:
        begin
            RED=8'hA0;
            GRN=8'h4B;
            BLU=8'h4E;
        end
        2072:
        begin
            RED=8'hDE;
            GRN=8'hE3;
            BLU=8'hDF;
        end
        2073:
        begin
            RED=8'hEF;
            GRN=8'hEF;
            BLU=8'hC9;
        end
        2074:
        begin
            RED=8'h2B;
            GRN=8'h29;
            BLU=8'h2C;
        end
        2075:
        begin
            RED=8'h24;
            GRN=8'h24;
            BLU=8'h24;
        end
        2076:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h25;
        end
        2077:
        begin
            RED=8'h21;
            GRN=8'h21;
            BLU=8'h23;
        end
        2078:
        begin
            RED=8'h21;
            GRN=8'h21;
            BLU=8'h23;
        end
        2079:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h20;
        end
        2080:
        begin
            RED=8'h1F;
            GRN=8'h1F;
            BLU=8'h1F;
        end
        2081:
        begin
            RED=8'h1E;
            GRN=8'h1E;
            BLU=8'h1E;
        end
        2082:
        begin
            RED=8'h1E;
            GRN=8'h1E;
            BLU=8'h1E;
        end
        2083:
        begin
            RED=8'h11;
            GRN=8'h11;
            BLU=8'h11;
        end
        2084:
        begin
            RED=8'h14;
            GRN=8'h14;
            BLU=8'h14;
        end
        2085:
        begin
            RED=8'h12;
            GRN=8'h10;
            BLU=8'h25;
        end
        2086:
        begin
            RED=8'h10;
            GRN=8'h0E;
            BLU=8'h1B;
        end
        2087:
        begin
            RED=8'h0D;
            GRN=8'h0C;
            BLU=8'h14;
        end
        2112:
        begin
            RED=8'h15;
            GRN=8'h14;
            BLU=8'h19;
        end
        2113:
        begin
            RED=8'h19;
            GRN=8'h19;
            BLU=8'h19;
        end
        2114:
        begin
            RED=8'h1F;
            GRN=8'h1F;
            BLU=8'h1F;
        end
        2115:
        begin
            RED=8'h24;
            GRN=8'h24;
            BLU=8'h26;
        end
        2116:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2117:
        begin
            RED=8'h2B;
            GRN=8'h2B;
            BLU=8'h2B;
        end
        2118:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        2119:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2C;
        end
        2120:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2C;
        end
        2121:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        2122:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        2123:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        2124:
        begin
            RED=8'h2B;
            GRN=8'h2B;
            BLU=8'h2D;
        end
        2125:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2C;
        end
        2126:
        begin
            RED=8'h27;
            GRN=8'h27;
            BLU=8'h27;
        end
        2127:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h29;
        end
        2128:
        begin
            RED=8'h2D;
            GRN=8'h2D;
            BLU=8'h2D;
        end
        2129:
        begin
            RED=8'h2B;
            GRN=8'h2B;
            BLU=8'h2B;
        end
        2130:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2131:
        begin
            RED=8'h55;
            GRN=8'h53;
            BLU=8'h44;
        end
        2132:
        begin
            RED=8'hED;
            GRN=8'hEC;
            BLU=8'hEA;
        end
        2133:
        begin
            RED=8'hD1;
            GRN=8'hD1;
            BLU=8'hD1;
        end
        2134:
        begin
            RED=8'h3C;
            GRN=8'h2A;
            BLU=8'h36;
        end
        2135:
        begin
            RED=8'h5E;
            GRN=8'h34;
            BLU=8'h40;
        end
        2136:
        begin
            RED=8'hE1;
            GRN=8'hE5;
            BLU=8'hE4;
        end
        2137:
        begin
            RED=8'hF6;
            GRN=8'hF7;
            BLU=8'hF2;
        end
        2138:
        begin
            RED=8'h29;
            GRN=8'h25;
            BLU=8'h24;
        end
        2139:
        begin
            RED=8'h25;
            GRN=8'h25;
            BLU=8'h25;
        end
        2140:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h23;
        end
        2141:
        begin
            RED=8'h22;
            GRN=8'h22;
            BLU=8'h24;
        end
        2142:
        begin
            RED=8'h24;
            GRN=8'h24;
            BLU=8'h24;
        end
        2143:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h20;
        end
        2144:
        begin
            RED=8'h1E;
            GRN=8'h1E;
            BLU=8'h1E;
        end
        2145:
        begin
            RED=8'h1F;
            GRN=8'h1F;
            BLU=8'h1F;
        end
        2146:
        begin
            RED=8'h1D;
            GRN=8'h1D;
            BLU=8'h1D;
        end
        2147:
        begin
            RED=8'h14;
            GRN=8'h14;
            BLU=8'h14;
        end
        2148:
        begin
            RED=8'h17;
            GRN=8'h17;
            BLU=8'h17;
        end
        2149:
        begin
            RED=8'h12;
            GRN=8'h12;
            BLU=8'h1A;
        end
        2150:
        begin
            RED=8'h11;
            GRN=8'h0E;
            BLU=8'h1F;
        end
        2151:
        begin
            RED=8'h0F;
            GRN=8'h0D;
            BLU=8'h1A;
        end
        2176:
        begin
            RED=8'h15;
            GRN=8'h15;
            BLU=8'h15;
        end
        2177:
        begin
            RED=8'h1A;
            GRN=8'h1A;
            BLU=8'h1A;
        end
        2178:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h22;
        end
        2179:
        begin
            RED=8'h25;
            GRN=8'h25;
            BLU=8'h25;
        end
        2180:
        begin
            RED=8'h27;
            GRN=8'h27;
            BLU=8'h27;
        end
        2181:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        2182:
        begin
            RED=8'h2C;
            GRN=8'h2C;
            BLU=8'h2E;
        end
        2183:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        2184:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2C;
        end
        2185:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        2186:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2C;
        end
        2187:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2C;
        end
        2188:
        begin
            RED=8'h2B;
            GRN=8'h2B;
            BLU=8'h2D;
        end
        2189:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2C;
        end
        2190:
        begin
            RED=8'h27;
            GRN=8'h27;
            BLU=8'h27;
        end
        2191:
        begin
            RED=8'h27;
            GRN=8'h27;
            BLU=8'h27;
        end
        2192:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        2193:
        begin
            RED=8'h2B;
            GRN=8'h2B;
            BLU=8'h2B;
        end
        2194:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h29;
        end
        2195:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2196:
        begin
            RED=8'hF7;
            GRN=8'hF9;
            BLU=8'hF4;
        end
        2197:
        begin
            RED=8'hE6;
            GRN=8'hE7;
            BLU=8'hE1;
        end
        2198:
        begin
            RED=8'hA1;
            GRN=8'h4A;
            BLU=8'h39;
        end
        2199:
        begin
            RED=8'h9B;
            GRN=8'h4C;
            BLU=8'h45;
        end
        2200:
        begin
            RED=8'h32;
            GRN=8'h25;
            BLU=8'h2F;
        end
        2201:
        begin
            RED=8'hF7;
            GRN=8'hF7;
            BLU=8'hF5;
        end
        2202:
        begin
            RED=8'hF6;
            GRN=8'hF2;
            BLU=8'hEF;
        end
        2203:
        begin
            RED=8'h25;
            GRN=8'h25;
            BLU=8'h25;
        end
        2204:
        begin
            RED=8'h22;
            GRN=8'h22;
            BLU=8'h22;
        end
        2205:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h25;
        end
        2206:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h25;
        end
        2207:
        begin
            RED=8'h22;
            GRN=8'h22;
            BLU=8'h24;
        end
        2208:
        begin
            RED=8'h1D;
            GRN=8'h1D;
            BLU=8'h1D;
        end
        2209:
        begin
            RED=8'h1E;
            GRN=8'h1E;
            BLU=8'h1E;
        end
        2210:
        begin
            RED=8'h1D;
            GRN=8'h1D;
            BLU=8'h1D;
        end
        2211:
        begin
            RED=8'h13;
            GRN=8'h13;
            BLU=8'h13;
        end
        2212:
        begin
            RED=8'h15;
            GRN=8'h15;
            BLU=8'h15;
        end
        2213:
        begin
            RED=8'h12;
            GRN=8'h12;
            BLU=8'h12;
        end
        2214:
        begin
            RED=8'h0F;
            GRN=8'h0C;
            BLU=8'h1D;
        end
        2215:
        begin
            RED=8'h0E;
            GRN=8'h0C;
            BLU=8'h19;
        end
        2240:
        begin
            RED=8'h14;
            GRN=8'h14;
            BLU=8'h14;
        end
        2241:
        begin
            RED=8'h1D;
            GRN=8'h1D;
            BLU=8'h1D;
        end
        2242:
        begin
            RED=8'h21;
            GRN=8'h21;
            BLU=8'h23;
        end
        2243:
        begin
            RED=8'h25;
            GRN=8'h25;
            BLU=8'h25;
        end
        2244:
        begin
            RED=8'h25;
            GRN=8'h25;
            BLU=8'h25;
        end
        2245:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h29;
        end
        2246:
        begin
            RED=8'h2C;
            GRN=8'h2C;
            BLU=8'h2E;
        end
        2247:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2C;
        end
        2248:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        2249:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h29;
        end
        2250:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h2A;
        end
        2251:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2C;
        end
        2252:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2C;
        end
        2253:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        2254:
        begin
            RED=8'h1D;
            GRN=8'h1D;
            BLU=8'h1D;
        end
        2255:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2256:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2257:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2C;
        end
        2258:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2259:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2260:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2C;
        end
        2261:
        begin
            RED=8'hF0;
            GRN=8'hF1;
            BLU=8'hEB;
        end
        2262:
        begin
            RED=8'h9D;
            GRN=8'h49;
            BLU=8'h2D;
        end
        2263:
        begin
            RED=8'h5A;
            GRN=8'h1D;
            BLU=8'h22;
        end
        2264:
        begin
            RED=8'h54;
            GRN=8'h34;
            BLU=8'h41;
        end
        2265:
        begin
            RED=8'hF3;
            GRN=8'hF3;
            BLU=8'hF1;
        end
        2266:
        begin
            RED=8'hF2;
            GRN=8'hF3;
            BLU=8'hEE;
        end
        2267:
        begin
            RED=8'h26;
            GRN=8'h26;
            BLU=8'h26;
        end
        2268:
        begin
            RED=8'h25;
            GRN=8'h25;
            BLU=8'h25;
        end
        2269:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h25;
        end
        2270:
        begin
            RED=8'h21;
            GRN=8'h21;
            BLU=8'h23;
        end
        2271:
        begin
            RED=8'h21;
            GRN=8'h21;
            BLU=8'h23;
        end
        2272:
        begin
            RED=8'h1F;
            GRN=8'h1F;
            BLU=8'h1F;
        end
        2273:
        begin
            RED=8'h1D;
            GRN=8'h1D;
            BLU=8'h1D;
        end
        2274:
        begin
            RED=8'h1C;
            GRN=8'h1C;
            BLU=8'h1C;
        end
        2275:
        begin
            RED=8'h16;
            GRN=8'h16;
            BLU=8'h16;
        end
        2276:
        begin
            RED=8'h15;
            GRN=8'h15;
            BLU=8'h15;
        end
        2277:
        begin
            RED=8'h13;
            GRN=8'h13;
            BLU=8'h13;
        end
        2278:
        begin
            RED=8'h10;
            GRN=8'h0D;
            BLU=8'h1E;
        end
        2279:
        begin
            RED=8'h0E;
            GRN=8'h0C;
            BLU=8'h19;
        end
        2304:
        begin
            RED=8'h1A;
            GRN=8'h1A;
            BLU=8'h1A;
        end
        2305:
        begin
            RED=8'h1C;
            GRN=8'h1C;
            BLU=8'h1C;
        end
        2306:
        begin
            RED=8'h19;
            GRN=8'h19;
            BLU=8'h19;
        end
        2307:
        begin
            RED=8'h24;
            GRN=8'h24;
            BLU=8'h24;
        end
        2308:
        begin
            RED=8'h24;
            GRN=8'h24;
            BLU=8'h24;
        end
        2309:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2310:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2A;
        end
        2311:
        begin
            RED=8'h2D;
            GRN=8'h2D;
            BLU=8'h2B;
        end
        2312:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2A;
        end
        2313:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h29;
        end
        2314:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h29;
        end
        2315:
        begin
            RED=8'h27;
            GRN=8'h27;
            BLU=8'h27;
        end
        2316:
        begin
            RED=8'h2D;
            GRN=8'h2D;
            BLU=8'h2F;
        end
        2317:
        begin
            RED=8'h2B;
            GRN=8'h2B;
            BLU=8'h2D;
        end
        2318:
        begin
            RED=8'h26;
            GRN=8'h26;
            BLU=8'h26;
        end
        2319:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2320:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2A;
        end
        2321:
        begin
            RED=8'h25;
            GRN=8'h25;
            BLU=8'h25;
        end
        2322:
        begin
            RED=8'h25;
            GRN=8'h25;
            BLU=8'h25;
        end
        2323:
        begin
            RED=8'h26;
            GRN=8'h26;
            BLU=8'h26;
        end
        2324:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h29;
        end
        2325:
        begin
            RED=8'hC7;
            GRN=8'hCE;
            BLU=8'hC7;
        end
        2326:
        begin
            RED=8'hBD;
            GRN=8'h46;
            BLU=8'h30;
        end
        2327:
        begin
            RED=8'hAC;
            GRN=8'h51;
            BLU=8'h3E;
        end
        2328:
        begin
            RED=8'h46;
            GRN=8'h2E;
            BLU=8'h50;
        end
        2329:
        begin
            RED=8'hEC;
            GRN=8'hEF;
            BLU=8'hE8;
        end
        2330:
        begin
            RED=8'hFA;
            GRN=8'hFC;
            BLU=8'hF9;
        end
        2331:
        begin
            RED=8'h1E;
            GRN=8'h1E;
            BLU=8'h1E;
        end
        2332:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2333:
        begin
            RED=8'h22;
            GRN=8'h22;
            BLU=8'h22;
        end
        2334:
        begin
            RED=8'h22;
            GRN=8'h22;
            BLU=8'h24;
        end
        2335:
        begin
            RED=8'h24;
            GRN=8'h24;
            BLU=8'h26;
        end
        2336:
        begin
            RED=8'h1E;
            GRN=8'h1E;
            BLU=8'h1E;
        end
        2337:
        begin
            RED=8'h1C;
            GRN=8'h1C;
            BLU=8'h1C;
        end
        2338:
        begin
            RED=8'h1C;
            GRN=8'h1C;
            BLU=8'h1C;
        end
        2339:
        begin
            RED=8'h17;
            GRN=8'h17;
            BLU=8'h17;
        end
        2340:
        begin
            RED=8'h15;
            GRN=8'h15;
            BLU=8'h15;
        end
        2341:
        begin
            RED=8'h12;
            GRN=8'h12;
            BLU=8'h12;
        end
        2342:
        begin
            RED=8'h0F;
            GRN=8'h0D;
            BLU=8'h1B;
        end
        2343:
        begin
            RED=8'h0D;
            GRN=8'h0B;
            BLU=8'h18;
        end
        2368:
        begin
            RED=8'h16;
            GRN=8'h16;
            BLU=8'h16;
        end
        2369:
        begin
            RED=8'h1E;
            GRN=8'h1E;
            BLU=8'h1E;
        end
        2370:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h20;
        end
        2371:
        begin
            RED=8'h18;
            GRN=8'h18;
            BLU=8'h18;
        end
        2372:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h20;
        end
        2373:
        begin
            RED=8'h26;
            GRN=8'h26;
            BLU=8'h26;
        end
        2374:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h29;
        end
        2375:
        begin
            RED=8'h2B;
            GRN=8'h2B;
            BLU=8'h2B;
        end
        2376:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h29;
        end
        2377:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h29;
        end
        2378:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2A;
        end
        2379:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h2B;
        end
        2380:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2381:
        begin
            RED=8'h27;
            GRN=8'h27;
            BLU=8'h27;
        end
        2382:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2C;
        end
        2383:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2384:
        begin
            RED=8'h26;
            GRN=8'h26;
            BLU=8'h26;
        end
        2385:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2A;
        end
        2386:
        begin
            RED=8'h27;
            GRN=8'h27;
            BLU=8'h27;
        end
        2387:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2388:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2389:
        begin
            RED=8'h28;
            GRN=8'h2A;
            BLU=8'h29;
        end
        2390:
        begin
            RED=8'h4C;
            GRN=8'h21;
            BLU=8'h28;
        end
        2391:
        begin
            RED=8'h9C;
            GRN=8'h4E;
            BLU=8'h3A;
        end
        2392:
        begin
            RED=8'h6A;
            GRN=8'h33;
            BLU=8'h30;
        end
        2393:
        begin
            RED=8'h4A;
            GRN=8'h34;
            BLU=8'h40;
        end
        2394:
        begin
            RED=8'hFF;
            GRN=8'hFE;
            BLU=8'hFC;
        end
        2395:
        begin
            RED=8'h2B;
            GRN=8'h29;
            BLU=8'h2A;
        end
        2396:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h23;
        end
        2397:
        begin
            RED=8'h22;
            GRN=8'h22;
            BLU=8'h24;
        end
        2398:
        begin
            RED=8'h21;
            GRN=8'h21;
            BLU=8'h23;
        end
        2399:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h22;
        end
        2400:
        begin
            RED=8'h1C;
            GRN=8'h1C;
            BLU=8'h1C;
        end
        2401:
        begin
            RED=8'h1B;
            GRN=8'h1B;
            BLU=8'h1B;
        end
        2402:
        begin
            RED=8'h1C;
            GRN=8'h1C;
            BLU=8'h1C;
        end
        2403:
        begin
            RED=8'h18;
            GRN=8'h18;
            BLU=8'h18;
        end
        2404:
        begin
            RED=8'h14;
            GRN=8'h14;
            BLU=8'h14;
        end
        2405:
        begin
            RED=8'h12;
            GRN=8'h12;
            BLU=8'h12;
        end
        2406:
        begin
            RED=8'h0F;
            GRN=8'h0D;
            BLU=8'h18;
        end
        2407:
        begin
            RED=8'h0D;
            GRN=8'h0B;
            BLU=8'h18;
        end
        2432:
        begin
            RED=8'h13;
            GRN=8'h13;
            BLU=8'h13;
        end
        2433:
        begin
            RED=8'h19;
            GRN=8'h19;
            BLU=8'h19;
        end
        2434:
        begin
            RED=8'h1F;
            GRN=8'h1F;
            BLU=8'h1F;
        end
        2435:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h20;
        end
        2436:
        begin
            RED=8'h1B;
            GRN=8'h1B;
            BLU=8'h1B;
        end
        2437:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h23;
        end
        2438:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2439:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2A;
        end
        2440:
        begin
            RED=8'h2C;
            GRN=8'h2C;
            BLU=8'h2E;
        end
        2441:
        begin
            RED=8'h2B;
            GRN=8'h2B;
            BLU=8'h2D;
        end
        2442:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2C;
        end
        2443:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2444:
        begin
            RED=8'h27;
            GRN=8'h27;
            BLU=8'h27;
        end
        2445:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2446:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h29;
        end
        2447:
        begin
            RED=8'h26;
            GRN=8'h26;
            BLU=8'h26;
        end
        2448:
        begin
            RED=8'h26;
            GRN=8'h26;
            BLU=8'h26;
        end
        2449:
        begin
            RED=8'h27;
            GRN=8'h27;
            BLU=8'h27;
        end
        2450:
        begin
            RED=8'h26;
            GRN=8'h26;
            BLU=8'h26;
        end
        2451:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2452:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2453:
        begin
            RED=8'h26;
            GRN=8'h26;
            BLU=8'h26;
        end
        2454:
        begin
            RED=8'h1F;
            GRN=8'h28;
            BLU=8'h27;
        end
        2455:
        begin
            RED=8'h68;
            GRN=8'h3A;
            BLU=8'h54;
        end
        2456:
        begin
            RED=8'h71;
            GRN=8'h3B;
            BLU=8'h39;
        end
        2457:
        begin
            RED=8'h5A;
            GRN=8'h2E;
            BLU=8'h3D;
        end
        2458:
        begin
            RED=8'hFF;
            GRN=8'hFF;
            BLU=8'hFF;
        end
        2459:
        begin
            RED=8'h7C;
            GRN=8'h7D;
            BLU=8'h78;
        end
        2460:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h23;
        end
        2461:
        begin
            RED=8'h24;
            GRN=8'h24;
            BLU=8'h24;
        end
        2462:
        begin
            RED=8'h22;
            GRN=8'h22;
            BLU=8'h24;
        end
        2463:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h22;
        end
        2464:
        begin
            RED=8'h1C;
            GRN=8'h1C;
            BLU=8'h1C;
        end
        2465:
        begin
            RED=8'h1C;
            GRN=8'h1C;
            BLU=8'h1C;
        end
        2466:
        begin
            RED=8'h19;
            GRN=8'h19;
            BLU=8'h19;
        end
        2467:
        begin
            RED=8'h18;
            GRN=8'h18;
            BLU=8'h18;
        end
        2468:
        begin
            RED=8'h13;
            GRN=8'h13;
            BLU=8'h13;
        end
        2469:
        begin
            RED=8'h11;
            GRN=8'h11;
            BLU=8'h11;
        end
        2470:
        begin
            RED=8'h10;
            GRN=8'h10;
            BLU=8'h10;
        end
        2471:
        begin
            RED=8'h0C;
            GRN=8'h0A;
            BLU=8'h17;
        end
        2496:
        begin
            RED=8'h12;
            GRN=8'h12;
            BLU=8'h12;
        end
        2497:
        begin
            RED=8'h17;
            GRN=8'h17;
            BLU=8'h17;
        end
        2498:
        begin
            RED=8'h1D;
            GRN=8'h1D;
            BLU=8'h1D;
        end
        2499:
        begin
            RED=8'h1F;
            GRN=8'h1F;
            BLU=8'h1F;
        end
        2500:
        begin
            RED=8'h21;
            GRN=8'h21;
            BLU=8'h21;
        end
        2501:
        begin
            RED=8'h1B;
            GRN=8'h1B;
            BLU=8'h1B;
        end
        2502:
        begin
            RED=8'h26;
            GRN=8'h26;
            BLU=8'h26;
        end
        2503:
        begin
            RED=8'h27;
            GRN=8'h27;
            BLU=8'h27;
        end
        2504:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2505:
        begin
            RED=8'h2B;
            GRN=8'h2B;
            BLU=8'h2D;
        end
        2506:
        begin
            RED=8'h2A;
            GRN=8'h2A;
            BLU=8'h2C;
        end
        2507:
        begin
            RED=8'h27;
            GRN=8'h27;
            BLU=8'h27;
        end
        2508:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h29;
        end
        2509:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2510:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2511:
        begin
            RED=8'h26;
            GRN=8'h26;
            BLU=8'h26;
        end
        2512:
        begin
            RED=8'h22;
            GRN=8'h22;
            BLU=8'h22;
        end
        2513:
        begin
            RED=8'h25;
            GRN=8'h25;
            BLU=8'h25;
        end
        2514:
        begin
            RED=8'h27;
            GRN=8'h27;
            BLU=8'h27;
        end
        2515:
        begin
            RED=8'h29;
            GRN=8'h29;
            BLU=8'h29;
        end
        2516:
        begin
            RED=8'h28;
            GRN=8'h28;
            BLU=8'h28;
        end
        2517:
        begin
            RED=8'h26;
            GRN=8'h26;
            BLU=8'h26;
        end
        2518:
        begin
            RED=8'h29;
            GRN=8'h27;
            BLU=8'h28;
        end
        2519:
        begin
            RED=8'hA4;
            GRN=8'h50;
            BLU=8'h38;
        end
        2520:
        begin
            RED=8'h7E;
            GRN=8'h40;
            BLU=8'h33;
        end
        2521:
        begin
            RED=8'h4F;
            GRN=8'h3D;
            BLU=8'h53;
        end
        2522:
        begin
            RED=8'h51;
            GRN=8'h31;
            BLU=8'h3E;
        end
        2523:
        begin
            RED=8'hEE;
            GRN=8'hEE;
            BLU=8'hEC;
        end
        2524:
        begin
            RED=8'h26;
            GRN=8'h26;
            BLU=8'h26;
        end
        2525:
        begin
            RED=8'h24;
            GRN=8'h24;
            BLU=8'h24;
        end
        2526:
        begin
            RED=8'h23;
            GRN=8'h23;
            BLU=8'h25;
        end
        2527:
        begin
            RED=8'h20;
            GRN=8'h20;
            BLU=8'h20;
        end
        2528:
        begin
            RED=8'h1D;
            GRN=8'h1D;
            BLU=8'h1D;
        end
        2529:
        begin
            RED=8'h1A;
            GRN=8'h1A;
            BLU=8'h1A;
        end
        2530:
        begin
            RED=8'h1A;
            GRN=8'h1A;
            BLU=8'h1A;
        end
        2531:
        begin
            RED=8'h17;
            GRN=8'h17;
            BLU=8'h17;
        end
        2532:
        begin
            RED=8'h14;
            GRN=8'h14;
            BLU=8'h14;
        end
        2533:
        begin
            RED=8'h10;
            GRN=8'h10;
            BLU=8'h10;
        end
        2534:
        begin
            RED=8'h0F;
            GRN=8'h0F;
            BLU=8'h0D;
        end
        2535:
        begin
            RED=8'h0B;
            GRN=8'h09;
            BLU=8'h14;
        end
        default:
        begin
            RED=8'h00;
            GRN=8'h00;
            BLU=8'h00;
        end
    endcase
endmodule
