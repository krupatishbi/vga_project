module professor_farnsworth_64x64_rom(
    input  [5:0] x_idx,
    input  [5:0] y_idx,
    output reg [7:0] RED,
    output reg [7:0] GRN,
    output reg [7:0] BLU);
always @ (*)
    case ({y_idx,x_idx})
        0:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        3:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        4:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        5:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        6:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        7:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        8:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        9:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        10:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        11:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        12:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        13:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        14:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        15:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        16:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        17:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        18:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        19:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        20:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        21:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        22:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        23:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        24:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        25:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        26:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        27:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        28:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        29:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        30:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        31:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        32:
        begin
            RED=8'h7F;
            GRN=8'h82;
            BLU=8'h65;
        end
        33:
        begin
            RED=8'h7F;
            GRN=8'h82;
            BLU=8'h65;
        end
        34:
        begin
            RED=8'h80;
            GRN=8'h82;
            BLU=8'h64;
        end
        35:
        begin
            RED=8'h81;
            GRN=8'h82;
            BLU=8'h63;
        end
        36:
        begin
            RED=8'h81;
            GRN=8'h82;
            BLU=8'h61;
        end
        37:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h5C;
        end
        38:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h5E;
        end
        39:
        begin
            RED=8'h79;
            GRN=8'h83;
            BLU=8'h61;
        end
        40:
        begin
            RED=8'h79;
            GRN=8'h86;
            BLU=8'h65;
        end
        41:
        begin
            RED=8'h78;
            GRN=8'h84;
            BLU=8'h69;
        end
        42:
        begin
            RED=8'h7C;
            GRN=8'h83;
            BLU=8'h67;
        end
        43:
        begin
            RED=8'h81;
            GRN=8'h80;
            BLU=8'h62;
        end
        44:
        begin
            RED=8'h88;
            GRN=8'h80;
            BLU=8'h5E;
        end
        45:
        begin
            RED=8'h8F;
            GRN=8'h81;
            BLU=8'h5A;
        end
        46:
        begin
            RED=8'h93;
            GRN=8'h7F;
            BLU=8'h52;
        end
        47:
        begin
            RED=8'h93;
            GRN=8'h7F;
            BLU=8'h52;
        end
        48:
        begin
            RED=8'h95;
            GRN=8'h80;
            BLU=8'h53;
        end
        49:
        begin
            RED=8'h94;
            GRN=8'h7F;
            BLU=8'h52;
        end
        50:
        begin
            RED=8'h8E;
            GRN=8'h7F;
            BLU=8'h57;
        end
        51:
        begin
            RED=8'h87;
            GRN=8'h7F;
            BLU=8'h5B;
        end
        52:
        begin
            RED=8'h82;
            GRN=8'h81;
            BLU=8'h60;
        end
        53:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h67;
        end
        54:
        begin
            RED=8'h79;
            GRN=8'h83;
            BLU=8'h6A;
        end
        55:
        begin
            RED=8'h7A;
            GRN=8'h82;
            BLU=8'h6F;
        end
        56:
        begin
            RED=8'h7F;
            GRN=8'h84;
            BLU=8'h62;
        end
        57:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h5D;
        end
        58:
        begin
            RED=8'h46;
            GRN=8'h4C;
            BLU=8'h37;
        end
        59:
        begin
            RED=8'h2D;
            GRN=8'h30;
            BLU=8'h26;
        end
        60:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        61:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        62:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        63:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        64:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        65:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        66:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        67:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        68:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        69:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        70:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        71:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        72:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        73:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        74:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        75:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        76:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        77:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        78:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        79:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        80:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        81:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        82:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        83:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        84:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        85:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        86:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        87:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        88:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        89:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        90:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        91:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        92:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        93:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        94:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        95:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        96:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h64;
        end
        97:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h65;
        end
        98:
        begin
            RED=8'h7C;
            GRN=8'h84;
            BLU=8'h65;
        end
        99:
        begin
            RED=8'h7B;
            GRN=8'h84;
            BLU=8'h67;
        end
        100:
        begin
            RED=8'h7C;
            GRN=8'h84;
            BLU=8'h69;
        end
        101:
        begin
            RED=8'h7D;
            GRN=8'h81;
            BLU=8'h67;
        end
        102:
        begin
            RED=8'h82;
            GRN=8'h83;
            BLU=8'h65;
        end
        103:
        begin
            RED=8'h85;
            GRN=8'h80;
            BLU=8'h5E;
        end
        104:
        begin
            RED=8'h85;
            GRN=8'h7C;
            BLU=8'h56;
        end
        105:
        begin
            RED=8'h8F;
            GRN=8'h7F;
            BLU=8'h52;
        end
        106:
        begin
            RED=8'hAA;
            GRN=8'h95;
            BLU=8'h63;
        end
        107:
        begin
            RED=8'hC7;
            GRN=8'hAB;
            BLU=8'h77;
        end
        108:
        begin
            RED=8'hD9;
            GRN=8'hB7;
            BLU=8'h81;
        end
        109:
        begin
            RED=8'hE4;
            GRN=8'hBD;
            BLU=8'h85;
        end
        110:
        begin
            RED=8'hE7;
            GRN=8'hBF;
            BLU=8'h82;
        end
        111:
        begin
            RED=8'hE7;
            GRN=8'hBF;
            BLU=8'h82;
        end
        112:
        begin
            RED=8'hEB;
            GRN=8'hC3;
            BLU=8'h85;
        end
        113:
        begin
            RED=8'hE9;
            GRN=8'hC2;
            BLU=8'h84;
        end
        114:
        begin
            RED=8'hE7;
            GRN=8'hC0;
            BLU=8'h85;
        end
        115:
        begin
            RED=8'hDD;
            GRN=8'hBB;
            BLU=8'h82;
        end
        116:
        begin
            RED=8'hD0;
            GRN=8'hB5;
            BLU=8'h7E;
        end
        117:
        begin
            RED=8'hB6;
            GRN=8'hA0;
            BLU=8'h6C;
        end
        118:
        begin
            RED=8'h98;
            GRN=8'h87;
            BLU=8'h56;
        end
        119:
        begin
            RED=8'h87;
            GRN=8'h7D;
            BLU=8'h5B;
        end
        120:
        begin
            RED=8'h80;
            GRN=8'h83;
            BLU=8'h61;
        end
        121:
        begin
            RED=8'h79;
            GRN=8'h84;
            BLU=8'h68;
        end
        122:
        begin
            RED=8'h46;
            GRN=8'h4D;
            BLU=8'h3D;
        end
        123:
        begin
            RED=8'h2E;
            GRN=8'h30;
            BLU=8'h27;
        end
        124:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        125:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        126:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        127:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        128:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        129:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        130:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        131:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        132:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        133:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        134:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        135:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        136:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        137:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        138:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        139:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        140:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        141:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        142:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        143:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        144:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        145:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        146:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        147:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        148:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        149:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        150:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        151:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        152:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        153:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        154:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        155:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        156:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        157:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        158:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        159:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        160:
        begin
            RED=8'h7B;
            GRN=8'h84;
            BLU=8'h62;
        end
        161:
        begin
            RED=8'h7A;
            GRN=8'h84;
            BLU=8'h62;
        end
        162:
        begin
            RED=8'h7B;
            GRN=8'h84;
            BLU=8'h63;
        end
        163:
        begin
            RED=8'h7A;
            GRN=8'h83;
            BLU=8'h62;
        end
        164:
        begin
            RED=8'h7E;
            GRN=8'h84;
            BLU=8'h62;
        end
        165:
        begin
            RED=8'h81;
            GRN=8'h7D;
            BLU=8'h59;
        end
        166:
        begin
            RED=8'h9A;
            GRN=8'h8B;
            BLU=8'h5F;
        end
        167:
        begin
            RED=8'hC4;
            GRN=8'hAA;
            BLU=8'h75;
        end
        168:
        begin
            RED=8'hE0;
            GRN=8'hBC;
            BLU=8'h81;
        end
        169:
        begin
            RED=8'hE8;
            GRN=8'hC3;
            BLU=8'h83;
        end
        170:
        begin
            RED=8'hE9;
            GRN=8'hC1;
            BLU=8'h80;
        end
        171:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        172:
        begin
            RED=8'hF0;
            GRN=8'hBF;
            BLU=8'h7D;
        end
        173:
        begin
            RED=8'hF0;
            GRN=8'hBE;
            BLU=8'h7C;
        end
        174:
        begin
            RED=8'hF0;
            GRN=8'hC0;
            BLU=8'h7C;
        end
        175:
        begin
            RED=8'hF0;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        176:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h7C;
        end
        177:
        begin
            RED=8'hEE;
            GRN=8'hBE;
            BLU=8'h7B;
        end
        178:
        begin
            RED=8'hF0;
            GRN=8'hBF;
            BLU=8'h7A;
        end
        179:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h7A;
        end
        180:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7C;
        end
        181:
        begin
            RED=8'hE9;
            GRN=8'hC1;
            BLU=8'h7E;
        end
        182:
        begin
            RED=8'hE8;
            GRN=8'hC2;
            BLU=8'h81;
        end
        183:
        begin
            RED=8'hD3;
            GRN=8'hB2;
            BLU=8'h7C;
        end
        184:
        begin
            RED=8'h8C;
            GRN=8'h84;
            BLU=8'h59;
        end
        185:
        begin
            RED=8'h7B;
            GRN=8'h82;
            BLU=8'h67;
        end
        186:
        begin
            RED=8'h4A;
            GRN=8'h4E;
            BLU=8'h41;
        end
        187:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        188:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        189:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        190:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        191:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        192:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        193:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        194:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        195:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        196:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        197:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        198:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        199:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        200:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        201:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        202:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        203:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        204:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        205:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        206:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        207:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        208:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        209:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        210:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        211:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        212:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        213:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        214:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        215:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        216:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        217:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        218:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        219:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        220:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        221:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        222:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        223:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        224:
        begin
            RED=8'h7D;
            GRN=8'h85;
            BLU=8'h65;
        end
        225:
        begin
            RED=8'h80;
            GRN=8'h84;
            BLU=8'h62;
        end
        226:
        begin
            RED=8'h85;
            GRN=8'h81;
            BLU=8'h59;
        end
        227:
        begin
            RED=8'h8E;
            GRN=8'h83;
            BLU=8'h55;
        end
        228:
        begin
            RED=8'hAE;
            GRN=8'h9C;
            BLU=8'h69;
        end
        229:
        begin
            RED=8'hDB;
            GRN=8'hBE;
            BLU=8'h82;
        end
        230:
        begin
            RED=8'hE7;
            GRN=8'hC6;
            BLU=8'h87;
        end
        231:
        begin
            RED=8'hE9;
            GRN=8'hC2;
            BLU=8'h7E;
        end
        232:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h7A;
        end
        233:
        begin
            RED=8'hEB;
            GRN=8'hC2;
            BLU=8'h80;
        end
        234:
        begin
            RED=8'hEA;
            GRN=8'hC2;
            BLU=8'h83;
        end
        235:
        begin
            RED=8'hEB;
            GRN=8'hC2;
            BLU=8'h82;
        end
        236:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h82;
        end
        237:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h82;
        end
        238:
        begin
            RED=8'hEB;
            GRN=8'hC1;
            BLU=8'h81;
        end
        239:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h81;
        end
        240:
        begin
            RED=8'hEB;
            GRN=8'hC1;
            BLU=8'h81;
        end
        241:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h81;
        end
        242:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        243:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        244:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h7F;
        end
        245:
        begin
            RED=8'hE9;
            GRN=8'hC2;
            BLU=8'h7E;
        end
        246:
        begin
            RED=8'hE9;
            GRN=8'hC2;
            BLU=8'h7F;
        end
        247:
        begin
            RED=8'hEB;
            GRN=8'hBF;
            BLU=8'h80;
        end
        248:
        begin
            RED=8'hE4;
            GRN=8'hC2;
            BLU=8'h84;
        end
        249:
        begin
            RED=8'hAB;
            GRN=8'h99;
            BLU=8'h6D;
        end
        250:
        begin
            RED=8'h4F;
            GRN=8'h48;
            BLU=8'h38;
        end
        251:
        begin
            RED=8'h30;
            GRN=8'h2F;
            BLU=8'h29;
        end
        252:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        253:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        254:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        255:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        256:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        257:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        258:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        259:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        260:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        261:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        262:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        263:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        264:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        265:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        266:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        267:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        268:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        269:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        270:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        271:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        272:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        273:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        274:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        275:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        276:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        277:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        278:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        279:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        280:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        281:
        begin
            RED=8'h7F;
            GRN=8'h82;
            BLU=8'h64;
        end
        282:
        begin
            RED=8'h7F;
            GRN=8'h82;
            BLU=8'h64;
        end
        283:
        begin
            RED=8'h7F;
            GRN=8'h82;
            BLU=8'h63;
        end
        284:
        begin
            RED=8'h7E;
            GRN=8'h84;
            BLU=8'h64;
        end
        285:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h64;
        end
        286:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h63;
        end
        287:
        begin
            RED=8'h7F;
            GRN=8'h84;
            BLU=8'h61;
        end
        288:
        begin
            RED=8'h80;
            GRN=8'h80;
            BLU=8'h5E;
        end
        289:
        begin
            RED=8'h88;
            GRN=8'h7E;
            BLU=8'h58;
        end
        290:
        begin
            RED=8'hBF;
            GRN=8'hA9;
            BLU=8'h79;
        end
        291:
        begin
            RED=8'hE2;
            GRN=8'hBF;
            BLU=8'h86;
        end
        292:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h83;
        end
        293:
        begin
            RED=8'hF1;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        294:
        begin
            RED=8'hEE;
            GRN=8'hBE;
            BLU=8'h7F;
        end
        295:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h83;
        end
        296:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h84;
        end
        297:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h7F;
        end
        298:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h7F;
        end
        299:
        begin
            RED=8'hEE;
            GRN=8'hC1;
            BLU=8'h7F;
        end
        300:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h80;
        end
        301:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h80;
        end
        302:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        303:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        304:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        305:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        306:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        307:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        308:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        309:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h7C;
        end
        310:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        311:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        312:
        begin
            RED=8'hF4;
            GRN=8'hBF;
            BLU=8'h75;
        end
        313:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h82;
        end
        314:
        begin
            RED=8'h8D;
            GRN=8'h79;
            BLU=8'h60;
        end
        315:
        begin
            RED=8'h31;
            GRN=8'h2E;
            BLU=8'h27;
        end
        316:
        begin
            RED=8'h2F;
            GRN=8'h31;
            BLU=8'h29;
        end
        317:
        begin
            RED=8'h2F;
            GRN=8'h32;
            BLU=8'h29;
        end
        318:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        319:
        begin
            RED=8'h31;
            GRN=8'h31;
            BLU=8'h29;
        end
        320:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        321:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        322:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        323:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        324:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        325:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        326:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        327:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        328:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        329:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        330:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        331:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        332:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        333:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        334:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        335:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        336:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        337:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        338:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        339:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        340:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        341:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        342:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        343:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        344:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h65;
        end
        345:
        begin
            RED=8'h7F;
            GRN=8'h82;
            BLU=8'h66;
        end
        346:
        begin
            RED=8'h80;
            GRN=8'h81;
            BLU=8'h67;
        end
        347:
        begin
            RED=8'h81;
            GRN=8'h82;
            BLU=8'h66;
        end
        348:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        349:
        begin
            RED=8'h7A;
            GRN=8'h82;
            BLU=8'h63;
        end
        350:
        begin
            RED=8'h7C;
            GRN=8'h80;
            BLU=8'h59;
        end
        351:
        begin
            RED=8'h88;
            GRN=8'h82;
            BLU=8'h51;
        end
        352:
        begin
            RED=8'hBC;
            GRN=8'hA4;
            BLU=8'h6D;
        end
        353:
        begin
            RED=8'hE4;
            GRN=8'hC3;
            BLU=8'h8A;
        end
        354:
        begin
            RED=8'hE9;
            GRN=8'hC1;
            BLU=8'h84;
        end
        355:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        356:
        begin
            RED=8'hF0;
            GRN=8'hBF;
            BLU=8'h7D;
        end
        357:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        358:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        359:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        360:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        361:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        362:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        363:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        364:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        365:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        366:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        367:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        368:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        369:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        370:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        371:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        372:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        373:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        374:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h80;
        end
        375:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h82;
        end
        376:
        begin
            RED=8'hF2;
            GRN=8'hBE;
            BLU=8'h7B;
        end
        377:
        begin
            RED=8'hF0;
            GRN=8'hC0;
            BLU=8'h82;
        end
        378:
        begin
            RED=8'hDE;
            GRN=8'hBD;
            BLU=8'h8D;
        end
        379:
        begin
            RED=8'h4B;
            GRN=8'h41;
            BLU=8'h2E;
        end
        380:
        begin
            RED=8'h2F;
            GRN=8'h31;
            BLU=8'h2C;
        end
        381:
        begin
            RED=8'h2D;
            GRN=8'h34;
            BLU=8'h29;
        end
        382:
        begin
            RED=8'h2F;
            GRN=8'h32;
            BLU=8'h28;
        end
        383:
        begin
            RED=8'h33;
            GRN=8'h30;
            BLU=8'h29;
        end
        384:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        385:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        386:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        387:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        388:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        389:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        390:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        391:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        392:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        393:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        394:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        395:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        396:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        397:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        398:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        399:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        400:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        401:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        402:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        403:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        404:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        405:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        406:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        407:
        begin
            RED=8'h7F;
            GRN=8'h82;
            BLU=8'h65;
        end
        408:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h65;
        end
        409:
        begin
            RED=8'h7C;
            GRN=8'h84;
            BLU=8'h64;
        end
        410:
        begin
            RED=8'h7B;
            GRN=8'h85;
            BLU=8'h64;
        end
        411:
        begin
            RED=8'h7C;
            GRN=8'h83;
            BLU=8'h64;
        end
        412:
        begin
            RED=8'h84;
            GRN=8'h84;
            BLU=8'h67;
        end
        413:
        begin
            RED=8'h82;
            GRN=8'h7A;
            BLU=8'h54;
        end
        414:
        begin
            RED=8'hB1;
            GRN=8'h9A;
            BLU=8'h67;
        end
        415:
        begin
            RED=8'hE0;
            GRN=8'hBD;
            BLU=8'h81;
        end
        416:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h87;
        end
        417:
        begin
            RED=8'hED;
            GRN=8'hBE;
            BLU=8'h85;
        end
        418:
        begin
            RED=8'hEE;
            GRN=8'hBE;
            BLU=8'h82;
        end
        419:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        420:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        421:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        422:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        423:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        424:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        425:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        426:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        427:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        428:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        429:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        430:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        431:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        432:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        433:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        434:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        435:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        436:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        437:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        438:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        439:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h83;
        end
        440:
        begin
            RED=8'hF0;
            GRN=8'hBF;
            BLU=8'h7C;
        end
        441:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7B;
        end
        442:
        begin
            RED=8'hE8;
            GRN=8'hC3;
            BLU=8'h84;
        end
        443:
        begin
            RED=8'h7F;
            GRN=8'h70;
            BLU=8'h51;
        end
        444:
        begin
            RED=8'h2F;
            GRN=8'h2E;
            BLU=8'h25;
        end
        445:
        begin
            RED=8'h2E;
            GRN=8'h32;
            BLU=8'h2A;
        end
        446:
        begin
            RED=8'h2F;
            GRN=8'h32;
            BLU=8'h2A;
        end
        447:
        begin
            RED=8'h32;
            GRN=8'h30;
            BLU=8'h28;
        end
        448:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        449:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        450:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        451:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        452:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        453:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        454:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        455:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        456:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        457:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        458:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        459:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        460:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        461:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        462:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        463:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        464:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        465:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        466:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        467:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        468:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        469:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        470:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        471:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h67;
        end
        472:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h65;
        end
        473:
        begin
            RED=8'h7D;
            GRN=8'h82;
            BLU=8'h60;
        end
        474:
        begin
            RED=8'h82;
            GRN=8'h88;
            BLU=8'h63;
        end
        475:
        begin
            RED=8'h81;
            GRN=8'h81;
            BLU=8'h5C;
        end
        476:
        begin
            RED=8'h8D;
            GRN=8'h7E;
            BLU=8'h56;
        end
        477:
        begin
            RED=8'hD2;
            GRN=8'hB4;
            BLU=8'h82;
        end
        478:
        begin
            RED=8'hEB;
            GRN=8'hBF;
            BLU=8'h82;
        end
        479:
        begin
            RED=8'hF2;
            GRN=8'hBE;
            BLU=8'h7C;
        end
        480:
        begin
            RED=8'hF2;
            GRN=8'hBD;
            BLU=8'h80;
        end
        481:
        begin
            RED=8'hF2;
            GRN=8'hBD;
            BLU=8'h82;
        end
        482:
        begin
            RED=8'hF0;
            GRN=8'hBE;
            BLU=8'h81;
        end
        483:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        484:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        485:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        486:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        487:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        488:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        489:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        490:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        491:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        492:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        493:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        494:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        495:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        496:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        497:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        498:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        499:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        500:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        501:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        502:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        503:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h82;
        end
        504:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        505:
        begin
            RED=8'hEF;
            GRN=8'hC0;
            BLU=8'h7B;
        end
        506:
        begin
            RED=8'hEC;
            GRN=8'hC2;
            BLU=8'h7B;
        end
        507:
        begin
            RED=8'hAC;
            GRN=8'h97;
            BLU=8'h6F;
        end
        508:
        begin
            RED=8'h31;
            GRN=8'h2C;
            BLU=8'h1F;
        end
        509:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h2B;
        end
        510:
        begin
            RED=8'h2F;
            GRN=8'h31;
            BLU=8'h2B;
        end
        511:
        begin
            RED=8'h31;
            GRN=8'h31;
            BLU=8'h27;
        end
        512:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        513:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        514:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        515:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        516:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        517:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        518:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        519:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        520:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        521:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        522:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        523:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        524:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        525:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        526:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        527:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        528:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        529:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        530:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        531:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        532:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        533:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        534:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        535:
        begin
            RED=8'h7C;
            GRN=8'h83;
            BLU=8'h68;
        end
        536:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h65;
        end
        537:
        begin
            RED=8'h84;
            GRN=8'h81;
            BLU=8'h60;
        end
        538:
        begin
            RED=8'h86;
            GRN=8'h7D;
            BLU=8'h59;
        end
        539:
        begin
            RED=8'hA7;
            GRN=8'h94;
            BLU=8'h65;
        end
        540:
        begin
            RED=8'hE2;
            GRN=8'hC2;
            BLU=8'h84;
        end
        541:
        begin
            RED=8'hEE;
            GRN=8'hC3;
            BLU=8'h81;
        end
        542:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h7D;
        end
        543:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        544:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        545:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        546:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        547:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h80;
        end
        548:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h80;
        end
        549:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        550:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        551:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        552:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        553:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        554:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        555:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        556:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        557:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        558:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        559:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        560:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        561:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        562:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        563:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        564:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        565:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        566:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        567:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h7F;
        end
        568:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        569:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        570:
        begin
            RED=8'hF0;
            GRN=8'hBE;
            BLU=8'h81;
        end
        571:
        begin
            RED=8'hB9;
            GRN=8'h9D;
            BLU=8'h75;
        end
        572:
        begin
            RED=8'h39;
            GRN=8'h31;
            BLU=8'h21;
        end
        573:
        begin
            RED=8'h31;
            GRN=8'h2F;
            BLU=8'h2B;
        end
        574:
        begin
            RED=8'h2F;
            GRN=8'h31;
            BLU=8'h2C;
        end
        575:
        begin
            RED=8'h31;
            GRN=8'h31;
            BLU=8'h26;
        end
        576:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        577:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        578:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        579:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        580:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        581:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        582:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        583:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        584:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        585:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        586:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        587:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        588:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        589:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        590:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        591:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        592:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        593:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        594:
        begin
            RED=8'h81;
            GRN=8'h82;
            BLU=8'h60;
        end
        595:
        begin
            RED=8'h81;
            GRN=8'h82;
            BLU=8'h61;
        end
        596:
        begin
            RED=8'h7D;
            GRN=8'h83;
            BLU=8'h67;
        end
        597:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h66;
        end
        598:
        begin
            RED=8'h81;
            GRN=8'h82;
            BLU=8'h62;
        end
        599:
        begin
            RED=8'h7F;
            GRN=8'h85;
            BLU=8'h6E;
        end
        600:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h63;
        end
        601:
        begin
            RED=8'h83;
            GRN=8'h7C;
            BLU=8'h50;
        end
        602:
        begin
            RED=8'hC5;
            GRN=8'hA5;
            BLU=8'h73;
        end
        603:
        begin
            RED=8'hEB;
            GRN=8'hC0;
            BLU=8'h86;
        end
        604:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h7E;
        end
        605:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7C;
        end
        606:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        607:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h81;
        end
        608:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        609:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        610:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        611:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        612:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        613:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        614:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        615:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        616:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        617:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        618:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        619:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        620:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        621:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        622:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        623:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        624:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        625:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        626:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        627:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        628:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        629:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        630:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        631:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h7D;
        end
        632:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h86;
        end
        633:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h80;
        end
        634:
        begin
            RED=8'hEC;
            GRN=8'hBE;
            BLU=8'h7F;
        end
        635:
        begin
            RED=8'hAE;
            GRN=8'h96;
            BLU=8'h73;
        end
        636:
        begin
            RED=8'h32;
            GRN=8'h2F;
            BLU=8'h1F;
        end
        637:
        begin
            RED=8'h2F;
            GRN=8'h2F;
            BLU=8'h26;
        end
        638:
        begin
            RED=8'h2F;
            GRN=8'h31;
            BLU=8'h2C;
        end
        639:
        begin
            RED=8'h2F;
            GRN=8'h31;
            BLU=8'h2B;
        end
        640:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        641:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        642:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        643:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        644:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        645:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        646:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        647:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        648:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        649:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        650:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        651:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        652:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        653:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        654:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        655:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        656:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        657:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        658:
        begin
            RED=8'h80;
            GRN=8'h82;
            BLU=8'h63;
        end
        659:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h65;
        end
        660:
        begin
            RED=8'h7B;
            GRN=8'h84;
            BLU=8'h6A;
        end
        661:
        begin
            RED=8'h7D;
            GRN=8'h83;
            BLU=8'h66;
        end
        662:
        begin
            RED=8'h81;
            GRN=8'h82;
            BLU=8'h61;
        end
        663:
        begin
            RED=8'h80;
            GRN=8'h81;
            BLU=8'h61;
        end
        664:
        begin
            RED=8'h86;
            GRN=8'h7D;
            BLU=8'h55;
        end
        665:
        begin
            RED=8'hCE;
            GRN=8'hB2;
            BLU=8'h80;
        end
        666:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h84;
        end
        667:
        begin
            RED=8'hEE;
            GRN=8'hBE;
            BLU=8'h7E;
        end
        668:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        669:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        670:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        671:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        672:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        673:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        674:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        675:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        676:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        677:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        678:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        679:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        680:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        681:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        682:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        683:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        684:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        685:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        686:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        687:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        688:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        689:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        690:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        691:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        692:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        693:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        694:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        695:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        696:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h86;
        end
        697:
        begin
            RED=8'hED;
            GRN=8'hC2;
            BLU=8'h80;
        end
        698:
        begin
            RED=8'hEA;
            GRN=8'hC0;
            BLU=8'h81;
        end
        699:
        begin
            RED=8'h90;
            GRN=8'h7E;
            BLU=8'h5E;
        end
        700:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h21;
        end
        701:
        begin
            RED=8'h30;
            GRN=8'h32;
            BLU=8'h26;
        end
        702:
        begin
            RED=8'h2F;
            GRN=8'h32;
            BLU=8'h2B;
        end
        703:
        begin
            RED=8'h2E;
            GRN=8'h32;
            BLU=8'h2D;
        end
        704:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        705:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        706:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        707:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        708:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        709:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        710:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        711:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        712:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        713:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        714:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        715:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        716:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        717:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        718:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        719:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        720:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        721:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        722:
        begin
            RED=8'h7D;
            GRN=8'h83;
            BLU=8'h66;
        end
        723:
        begin
            RED=8'h7C;
            GRN=8'h83;
            BLU=8'h67;
        end
        724:
        begin
            RED=8'h80;
            GRN=8'h82;
            BLU=8'h63;
        end
        725:
        begin
            RED=8'h7F;
            GRN=8'h7B;
            BLU=8'h56;
        end
        726:
        begin
            RED=8'h82;
            GRN=8'h7B;
            BLU=8'h53;
        end
        727:
        begin
            RED=8'h80;
            GRN=8'h75;
            BLU=8'h42;
        end
        728:
        begin
            RED=8'hC3;
            GRN=8'hA3;
            BLU=8'h70;
        end
        729:
        begin
            RED=8'hEE;
            GRN=8'hBD;
            BLU=8'h85;
        end
        730:
        begin
            RED=8'hED;
            GRN=8'hBE;
            BLU=8'h7D;
        end
        731:
        begin
            RED=8'hED;
            GRN=8'hC3;
            BLU=8'h7E;
        end
        732:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        733:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        734:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        735:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        736:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        737:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        738:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        739:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        740:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        741:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h82;
        end
        742:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h82;
        end
        743:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h81;
        end
        744:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h82;
        end
        745:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h7F;
        end
        746:
        begin
            RED=8'hEE;
            GRN=8'hC1;
            BLU=8'h80;
        end
        747:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        748:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        749:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        750:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        751:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        752:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        753:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        754:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        755:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        756:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        757:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        758:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        759:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        760:
        begin
            RED=8'hEF;
            GRN=8'hBE;
            BLU=8'h85;
        end
        761:
        begin
            RED=8'hEC;
            GRN=8'hC1;
            BLU=8'h7E;
        end
        762:
        begin
            RED=8'hE7;
            GRN=8'hC2;
            BLU=8'h87;
        end
        763:
        begin
            RED=8'h62;
            GRN=8'h53;
            BLU=8'h39;
        end
        764:
        begin
            RED=8'h30;
            GRN=8'h30;
            BLU=8'h23;
        end
        765:
        begin
            RED=8'h31;
            GRN=8'h33;
            BLU=8'h28;
        end
        766:
        begin
            RED=8'h2F;
            GRN=8'h32;
            BLU=8'h29;
        end
        767:
        begin
            RED=8'h2E;
            GRN=8'h32;
            BLU=8'h2A;
        end
        768:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        769:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        770:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        771:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        772:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        773:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        774:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        775:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        776:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        777:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        778:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        779:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        780:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        781:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        782:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        783:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        784:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        785:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        786:
        begin
            RED=8'h80;
            GRN=8'h84;
            BLU=8'h64;
        end
        787:
        begin
            RED=8'h83;
            GRN=8'h80;
            BLU=8'h5C;
        end
        788:
        begin
            RED=8'h94;
            GRN=8'h84;
            BLU=8'h55;
        end
        789:
        begin
            RED=8'hC7;
            GRN=8'hAF;
            BLU=8'h79;
        end
        790:
        begin
            RED=8'hDC;
            GRN=8'hC0;
            BLU=8'h89;
        end
        791:
        begin
            RED=8'hE3;
            GRN=8'hC1;
            BLU=8'h82;
        end
        792:
        begin
            RED=8'hE6;
            GRN=8'hBC;
            BLU=8'h7E;
        end
        793:
        begin
            RED=8'hEA;
            GRN=8'hB9;
            BLU=8'h7A;
        end
        794:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h7D;
        end
        795:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        796:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        797:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        798:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        799:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        800:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        801:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        802:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        803:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        804:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h80;
        end
        805:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h83;
        end
        806:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h83;
        end
        807:
        begin
            RED=8'hEC;
            GRN=8'hBE;
            BLU=8'h82;
        end
        808:
        begin
            RED=8'hEC;
            GRN=8'hBE;
            BLU=8'h82;
        end
        809:
        begin
            RED=8'hE9;
            GRN=8'hBC;
            BLU=8'h7D;
        end
        810:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        811:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        812:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        813:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        814:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        815:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        816:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        817:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        818:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        819:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        820:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        821:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        822:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        823:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        824:
        begin
            RED=8'hF0;
            GRN=8'hBE;
            BLU=8'h83;
        end
        825:
        begin
            RED=8'hEC;
            GRN=8'hBE;
            BLU=8'h7C;
        end
        826:
        begin
            RED=8'hDF;
            GRN=8'hC0;
            BLU=8'h89;
        end
        827:
        begin
            RED=8'h42;
            GRN=8'h36;
            BLU=8'h23;
        end
        828:
        begin
            RED=8'h30;
            GRN=8'h30;
            BLU=8'h26;
        end
        829:
        begin
            RED=8'h31;
            GRN=8'h32;
            BLU=8'h28;
        end
        830:
        begin
            RED=8'h2F;
            GRN=8'h32;
            BLU=8'h27;
        end
        831:
        begin
            RED=8'h2E;
            GRN=8'h33;
            BLU=8'h27;
        end
        832:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        833:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        834:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        835:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        836:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        837:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        838:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        839:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        840:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        841:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        842:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        843:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h62;
        end
        844:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h62;
        end
        845:
        begin
            RED=8'h7D;
            GRN=8'h83;
            BLU=8'h62;
        end
        846:
        begin
            RED=8'h7C;
            GRN=8'h84;
            BLU=8'h63;
        end
        847:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h65;
        end
        848:
        begin
            RED=8'h80;
            GRN=8'h82;
            BLU=8'h65;
        end
        849:
        begin
            RED=8'h7F;
            GRN=8'h81;
            BLU=8'h60;
        end
        850:
        begin
            RED=8'h7F;
            GRN=8'h7A;
            BLU=8'h54;
        end
        851:
        begin
            RED=8'hAE;
            GRN=8'h9A;
            BLU=8'h6A;
        end
        852:
        begin
            RED=8'hDF;
            GRN=8'hBC;
            BLU=8'h7F;
        end
        853:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h7F;
        end
        854:
        begin
            RED=8'hEF;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        855:
        begin
            RED=8'hF1;
            GRN=8'hBF;
            BLU=8'h7D;
        end
        856:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h7D;
        end
        857:
        begin
            RED=8'hE8;
            GRN=8'hC3;
            BLU=8'h7F;
        end
        858:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h81;
        end
        859:
        begin
            RED=8'hF0;
            GRN=8'hBE;
            BLU=8'h80;
        end
        860:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        861:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        862:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        863:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        864:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        865:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        866:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        867:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        868:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        869:
        begin
            RED=8'hEB;
            GRN=8'hBE;
            BLU=8'h82;
        end
        870:
        begin
            RED=8'hD8;
            GRN=8'hAB;
            BLU=8'h6F;
        end
        871:
        begin
            RED=8'hD6;
            GRN=8'hA9;
            BLU=8'h6D;
        end
        872:
        begin
            RED=8'hD8;
            GRN=8'hAA;
            BLU=8'h6F;
        end
        873:
        begin
            RED=8'hD7;
            GRN=8'hAA;
            BLU=8'h6A;
        end
        874:
        begin
            RED=8'hD5;
            GRN=8'hA8;
            BLU=8'h67;
        end
        875:
        begin
            RED=8'hEB;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        876:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        877:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        878:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        879:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        880:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        881:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        882:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        883:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        884:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        885:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        886:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        887:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h80;
        end
        888:
        begin
            RED=8'hF1;
            GRN=8'hBE;
            BLU=8'h80;
        end
        889:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h7E;
        end
        890:
        begin
            RED=8'hC6;
            GRN=8'hAD;
            BLU=8'h7D;
        end
        891:
        begin
            RED=8'h38;
            GRN=8'h30;
            BLU=8'h1F;
        end
        892:
        begin
            RED=8'h30;
            GRN=8'h30;
            BLU=8'h28;
        end
        893:
        begin
            RED=8'h31;
            GRN=8'h32;
            BLU=8'h28;
        end
        894:
        begin
            RED=8'h2F;
            GRN=8'h32;
            BLU=8'h26;
        end
        895:
        begin
            RED=8'h2E;
            GRN=8'h32;
            BLU=8'h26;
        end
        896:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        897:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        898:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        899:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        900:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        901:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        902:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        903:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        904:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        905:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h65;
        end
        906:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h63;
        end
        907:
        begin
            RED=8'h7E;
            GRN=8'h84;
            BLU=8'h60;
        end
        908:
        begin
            RED=8'h7E;
            GRN=8'h84;
            BLU=8'h60;
        end
        909:
        begin
            RED=8'h7C;
            GRN=8'h85;
            BLU=8'h60;
        end
        910:
        begin
            RED=8'h7A;
            GRN=8'h86;
            BLU=8'h61;
        end
        911:
        begin
            RED=8'h84;
            GRN=8'h7F;
            BLU=8'h68;
        end
        912:
        begin
            RED=8'h89;
            GRN=8'h74;
            BLU=8'h5B;
        end
        913:
        begin
            RED=8'hB1;
            GRN=8'h96;
            BLU=8'h67;
        end
        914:
        begin
            RED=8'hDA;
            GRN=8'hBA;
            BLU=8'h7B;
        end
        915:
        begin
            RED=8'hE2;
            GRN=8'hBA;
            BLU=8'h7B;
        end
        916:
        begin
            RED=8'hDE;
            GRN=8'hB5;
            BLU=8'h75;
        end
        917:
        begin
            RED=8'hD3;
            GRN=8'hAA;
            BLU=8'h6A;
        end
        918:
        begin
            RED=8'hEB;
            GRN=8'hC0;
            BLU=8'h80;
        end
        919:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        920:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        921:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        922:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        923:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        924:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        925:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        926:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        927:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        928:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        929:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        930:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        931:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        932:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h81;
        end
        933:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h80;
        end
        934:
        begin
            RED=8'hE9;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        935:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h7F;
        end
        936:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h7F;
        end
        937:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        938:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        939:
        begin
            RED=8'hE7;
            GRN=8'hBA;
            BLU=8'h79;
        end
        940:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        941:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        942:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        943:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        944:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        945:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        946:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        947:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        948:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        949:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        950:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h80;
        end
        951:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h81;
        end
        952:
        begin
            RED=8'hF0;
            GRN=8'hC0;
            BLU=8'h78;
        end
        953:
        begin
            RED=8'hE8;
            GRN=8'hC1;
            BLU=8'h84;
        end
        954:
        begin
            RED=8'h89;
            GRN=8'h7B;
            BLU=8'h5D;
        end
        955:
        begin
            RED=8'h31;
            GRN=8'h31;
            BLU=8'h25;
        end
        956:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        957:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        958:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        959:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        960:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        961:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        962:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        963:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        964:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        965:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        966:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        967:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        968:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        969:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h62;
        end
        970:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h62;
        end
        971:
        begin
            RED=8'h7B;
            GRN=8'h84;
            BLU=8'h65;
        end
        972:
        begin
            RED=8'h7B;
            GRN=8'h84;
            BLU=8'h67;
        end
        973:
        begin
            RED=8'h7B;
            GRN=8'h84;
            BLU=8'h65;
        end
        974:
        begin
            RED=8'h83;
            GRN=8'h7E;
            BLU=8'h5B;
        end
        975:
        begin
            RED=8'h96;
            GRN=8'h81;
            BLU=8'h53;
        end
        976:
        begin
            RED=8'hDF;
            GRN=8'hB8;
            BLU=8'h81;
        end
        977:
        begin
            RED=8'hEE;
            GRN=8'hBE;
            BLU=8'h80;
        end
        978:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h81;
        end
        979:
        begin
            RED=8'hEB;
            GRN=8'hBF;
            BLU=8'h80;
        end
        980:
        begin
            RED=8'hEE;
            GRN=8'hC3;
            BLU=8'h84;
        end
        981:
        begin
            RED=8'hEB;
            GRN=8'hC0;
            BLU=8'h81;
        end
        982:
        begin
            RED=8'hED;
            GRN=8'hC2;
            BLU=8'h82;
        end
        983:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        984:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        985:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        986:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        987:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        988:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        989:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        990:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        991:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        992:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        993:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        994:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        995:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        996:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h80;
        end
        997:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h80;
        end
        998:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h80;
        end
        999:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h80;
        end
        1000:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h80;
        end
        1001:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1002:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        1003:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1004:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1005:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1006:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1007:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1008:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1009:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1010:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1011:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1012:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1013:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1014:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h80;
        end
        1015:
        begin
            RED=8'hEB;
            GRN=8'hC1;
            BLU=8'h80;
        end
        1016:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h7C;
        end
        1017:
        begin
            RED=8'hE0;
            GRN=8'hBF;
            BLU=8'h86;
        end
        1018:
        begin
            RED=8'h54;
            GRN=8'h4A;
            BLU=8'h2F;
        end
        1019:
        begin
            RED=8'h30;
            GRN=8'h30;
            BLU=8'h27;
        end
        1020:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1021:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1022:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1023:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1024:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1025:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1026:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1027:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1028:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1029:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1030:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1031:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1032:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1033:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h5F;
        end
        1034:
        begin
            RED=8'h7C;
            GRN=8'h84;
            BLU=8'h63;
        end
        1035:
        begin
            RED=8'h79;
            GRN=8'h83;
            BLU=8'h68;
        end
        1036:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h66;
        end
        1037:
        begin
            RED=8'h83;
            GRN=8'h7F;
            BLU=8'h60;
        end
        1038:
        begin
            RED=8'h88;
            GRN=8'h7A;
            BLU=8'h59;
        end
        1039:
        begin
            RED=8'hD6;
            GRN=8'hBC;
            BLU=8'h88;
        end
        1040:
        begin
            RED=8'hE6;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        1041:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h82;
        end
        1042:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h83;
        end
        1043:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        1044:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        1045:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        1046:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h81;
        end
        1047:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1048:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1049:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1050:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1051:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1052:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1053:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1054:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1055:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1056:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h80;
        end
        1057:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h82;
        end
        1058:
        begin
            RED=8'hEA;
            GRN=8'hBC;
            BLU=8'h7E;
        end
        1059:
        begin
            RED=8'hD8;
            GRN=8'hAA;
            BLU=8'h6C;
        end
        1060:
        begin
            RED=8'hCB;
            GRN=8'h9F;
            BLU=8'h61;
        end
        1061:
        begin
            RED=8'hD1;
            GRN=8'hA8;
            BLU=8'h6A;
        end
        1062:
        begin
            RED=8'hD2;
            GRN=8'hA9;
            BLU=8'h6A;
        end
        1063:
        begin
            RED=8'hD5;
            GRN=8'hAC;
            BLU=8'h6E;
        end
        1064:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h82;
        end
        1065:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        1066:
        begin
            RED=8'hEE;
            GRN=8'hC1;
            BLU=8'h80;
        end
        1067:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1068:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1069:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1070:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1071:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1072:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1073:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1074:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1075:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1076:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1077:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1078:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1079:
        begin
            RED=8'hEC;
            GRN=8'hC1;
            BLU=8'h7F;
        end
        1080:
        begin
            RED=8'hEB;
            GRN=8'hC3;
            BLU=8'h82;
        end
        1081:
        begin
            RED=8'hCD;
            GRN=8'hB4;
            BLU=8'h83;
        end
        1082:
        begin
            RED=8'h4D;
            GRN=8'h49;
            BLU=8'h33;
        end
        1083:
        begin
            RED=8'h2E;
            GRN=8'h31;
            BLU=8'h28;
        end
        1084:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1085:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1086:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1087:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1088:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1089:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1090:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1091:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1092:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1093:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1094:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1095:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1096:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1097:
        begin
            RED=8'h7E;
            GRN=8'h84;
            BLU=8'h60;
        end
        1098:
        begin
            RED=8'h7B;
            GRN=8'h85;
            BLU=8'h64;
        end
        1099:
        begin
            RED=8'h7D;
            GRN=8'h83;
            BLU=8'h68;
        end
        1100:
        begin
            RED=8'h8B;
            GRN=8'h80;
            BLU=8'h5E;
        end
        1101:
        begin
            RED=8'hAF;
            GRN=8'h93;
            BLU=8'h66;
        end
        1102:
        begin
            RED=8'hCA;
            GRN=8'hAB;
            BLU=8'h7B;
        end
        1103:
        begin
            RED=8'hD7;
            GRN=8'hB0;
            BLU=8'h7B;
        end
        1104:
        begin
            RED=8'hD6;
            GRN=8'hAB;
            BLU=8'h6F;
        end
        1105:
        begin
            RED=8'hD4;
            GRN=8'hAC;
            BLU=8'h6C;
        end
        1106:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h80;
        end
        1107:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h81;
        end
        1108:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h81;
        end
        1109:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h81;
        end
        1110:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h81;
        end
        1111:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1112:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1113:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1114:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1115:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1116:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1117:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1118:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1119:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1120:
        begin
            RED=8'hEC;
            GRN=8'hBE;
            BLU=8'h80;
        end
        1121:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h82;
        end
        1122:
        begin
            RED=8'hD8;
            GRN=8'hAA;
            BLU=8'h6C;
        end
        1123:
        begin
            RED=8'hE7;
            GRN=8'hB9;
            BLU=8'h7B;
        end
        1124:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h81;
        end
        1125:
        begin
            RED=8'hEC;
            GRN=8'hC2;
            BLU=8'h86;
        end
        1126:
        begin
            RED=8'hEA;
            GRN=8'hC0;
            BLU=8'h84;
        end
        1127:
        begin
            RED=8'hE1;
            GRN=8'hB7;
            BLU=8'h7A;
        end
        1128:
        begin
            RED=8'hCC;
            GRN=8'hA2;
            BLU=8'h65;
        end
        1129:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h81;
        end
        1130:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1131:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1132:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1133:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1134:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1135:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1136:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1137:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1138:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1139:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1140:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1141:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1142:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        1143:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        1144:
        begin
            RED=8'hE7;
            GRN=8'hC4;
            BLU=8'h86;
        end
        1145:
        begin
            RED=8'h9F;
            GRN=8'h8D;
            BLU=8'h62;
        end
        1146:
        begin
            RED=8'h4F;
            GRN=8'h50;
            BLU=8'h3D;
        end
        1147:
        begin
            RED=8'h2F;
            GRN=8'h32;
            BLU=8'h2A;
        end
        1148:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1149:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1150:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1151:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1152:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1153:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1154:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1155:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1156:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        1157:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h66;
        end
        1158:
        begin
            RED=8'h7D;
            GRN=8'h85;
            BLU=8'h61;
        end
        1159:
        begin
            RED=8'h7D;
            GRN=8'h85;
            BLU=8'h61;
        end
        1160:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h65;
        end
        1161:
        begin
            RED=8'h7A;
            GRN=8'h84;
            BLU=8'h64;
        end
        1162:
        begin
            RED=8'h81;
            GRN=8'h83;
            BLU=8'h63;
        end
        1163:
        begin
            RED=8'h8D;
            GRN=8'h7D;
            BLU=8'h58;
        end
        1164:
        begin
            RED=8'hD7;
            GRN=8'hB7;
            BLU=8'h84;
        end
        1165:
        begin
            RED=8'hE8;
            GRN=8'hC1;
            BLU=8'h81;
        end
        1166:
        begin
            RED=8'hE8;
            GRN=8'hC2;
            BLU=8'h80;
        end
        1167:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h81;
        end
        1168:
        begin
            RED=8'hF1;
            GRN=8'hBE;
            BLU=8'h80;
        end
        1169:
        begin
            RED=8'hEC;
            GRN=8'hC1;
            BLU=8'h7C;
        end
        1170:
        begin
            RED=8'hE9;
            GRN=8'hC2;
            BLU=8'h7D;
        end
        1171:
        begin
            RED=8'hED;
            GRN=8'hC2;
            BLU=8'h80;
        end
        1172:
        begin
            RED=8'hEF;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1173:
        begin
            RED=8'hEC;
            GRN=8'hBE;
            BLU=8'h82;
        end
        1174:
        begin
            RED=8'hE4;
            GRN=8'hBA;
            BLU=8'h84;
        end
        1175:
        begin
            RED=8'hE9;
            GRN=8'hBE;
            BLU=8'h81;
        end
        1176:
        begin
            RED=8'hEA;
            GRN=8'hC2;
            BLU=8'h7F;
        end
        1177:
        begin
            RED=8'hEC;
            GRN=8'hC2;
            BLU=8'h7D;
        end
        1178:
        begin
            RED=8'hEE;
            GRN=8'hBE;
            BLU=8'h7F;
        end
        1179:
        begin
            RED=8'hF2;
            GRN=8'hBF;
            BLU=8'h84;
        end
        1180:
        begin
            RED=8'hEE;
            GRN=8'hBD;
            BLU=8'h80;
        end
        1181:
        begin
            RED=8'hED;
            GRN=8'hBE;
            BLU=8'h80;
        end
        1182:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h83;
        end
        1183:
        begin
            RED=8'hEC;
            GRN=8'hC1;
            BLU=8'h84;
        end
        1184:
        begin
            RED=8'hF0;
            GRN=8'hBE;
            BLU=8'h86;
        end
        1185:
        begin
            RED=8'hEB;
            GRN=8'hBF;
            BLU=8'h7F;
        end
        1186:
        begin
            RED=8'hE9;
            GRN=8'hC1;
            BLU=8'h7A;
        end
        1187:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7C;
        end
        1188:
        begin
            RED=8'hF1;
            GRN=8'hBF;
            BLU=8'h80;
        end
        1189:
        begin
            RED=8'hEB;
            GRN=8'hBF;
            BLU=8'h7F;
        end
        1190:
        begin
            RED=8'hE9;
            GRN=8'hC2;
            BLU=8'h7F;
        end
        1191:
        begin
            RED=8'hE8;
            GRN=8'hC2;
            BLU=8'h80;
        end
        1192:
        begin
            RED=8'hE1;
            GRN=8'hB7;
            BLU=8'h79;
        end
        1193:
        begin
            RED=8'hE6;
            GRN=8'hB9;
            BLU=8'h7A;
        end
        1194:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1195:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1196:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1197:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1198:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1199:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1200:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1201:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1202:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1203:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1204:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1205:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1206:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        1207:
        begin
            RED=8'hF0;
            GRN=8'hBF;
            BLU=8'h79;
        end
        1208:
        begin
            RED=8'hDE;
            GRN=8'hBF;
            BLU=8'h8A;
        end
        1209:
        begin
            RED=8'h81;
            GRN=8'h79;
            BLU=8'h53;
        end
        1210:
        begin
            RED=8'h50;
            GRN=8'h53;
            BLU=8'h42;
        end
        1211:
        begin
            RED=8'h2F;
            GRN=8'h31;
            BLU=8'h2B;
        end
        1212:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1213:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1214:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1215:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1216:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1217:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1218:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1219:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1220:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        1221:
        begin
            RED=8'h7F;
            GRN=8'h82;
            BLU=8'h65;
        end
        1222:
        begin
            RED=8'h7E;
            GRN=8'h84;
            BLU=8'h60;
        end
        1223:
        begin
            RED=8'h7E;
            GRN=8'h84;
            BLU=8'h60;
        end
        1224:
        begin
            RED=8'h7D;
            GRN=8'h83;
            BLU=8'h66;
        end
        1225:
        begin
            RED=8'h7B;
            GRN=8'h84;
            BLU=8'h66;
        end
        1226:
        begin
            RED=8'h83;
            GRN=8'h7C;
            BLU=8'h59;
        end
        1227:
        begin
            RED=8'hD5;
            GRN=8'hB6;
            BLU=8'h8A;
        end
        1228:
        begin
            RED=8'hEB;
            GRN=8'hC2;
            BLU=8'h88;
        end
        1229:
        begin
            RED=8'hEC;
            GRN=8'hC4;
            BLU=8'h7E;
        end
        1230:
        begin
            RED=8'hEF;
            GRN=8'hC0;
            BLU=8'h78;
        end
        1231:
        begin
            RED=8'hF1;
            GRN=8'hBE;
            BLU=8'h7C;
        end
        1232:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h7F;
        end
        1233:
        begin
            RED=8'hE8;
            GRN=8'hC1;
            BLU=8'h83;
        end
        1234:
        begin
            RED=8'hE7;
            GRN=8'hC2;
            BLU=8'h80;
        end
        1235:
        begin
            RED=8'hD1;
            GRN=8'hA9;
            BLU=8'h64;
        end
        1236:
        begin
            RED=8'hEB;
            GRN=8'hC2;
            BLU=8'h83;
        end
        1237:
        begin
            RED=8'hEA;
            GRN=8'hBE;
            BLU=8'h83;
        end
        1238:
        begin
            RED=8'hCD;
            GRN=8'hA0;
            BLU=8'h67;
        end
        1239:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7C;
        end
        1240:
        begin
            RED=8'hE4;
            GRN=8'hC3;
            BLU=8'h88;
        end
        1241:
        begin
            RED=8'hC8;
            GRN=8'hB6;
            BLU=8'h89;
        end
        1242:
        begin
            RED=8'hB5;
            GRN=8'hAA;
            BLU=8'h89;
        end
        1243:
        begin
            RED=8'hB3;
            GRN=8'hAA;
            BLU=8'h8D;
        end
        1244:
        begin
            RED=8'hB2;
            GRN=8'hA6;
            BLU=8'h89;
        end
        1245:
        begin
            RED=8'hBF;
            GRN=8'hAA;
            BLU=8'h84;
        end
        1246:
        begin
            RED=8'hD5;
            GRN=8'hB7;
            BLU=8'h85;
        end
        1247:
        begin
            RED=8'hE4;
            GRN=8'hBF;
            BLU=8'h85;
        end
        1248:
        begin
            RED=8'hF1;
            GRN=8'hC0;
            BLU=8'h83;
        end
        1249:
        begin
            RED=8'hEF;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        1250:
        begin
            RED=8'hEE;
            GRN=8'hC2;
            BLU=8'h7D;
        end
        1251:
        begin
            RED=8'hEC;
            GRN=8'hC1;
            BLU=8'h82;
        end
        1252:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h86;
        end
        1253:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h80;
        end
        1254:
        begin
            RED=8'hEA;
            GRN=8'hC5;
            BLU=8'h7E;
        end
        1255:
        begin
            RED=8'hE9;
            GRN=8'hC4;
            BLU=8'h7E;
        end
        1256:
        begin
            RED=8'hEB;
            GRN=8'hBF;
            BLU=8'h82;
        end
        1257:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h80;
        end
        1258:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1259:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1260:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1261:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1262:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1263:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1264:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1265:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1266:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1267:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1268:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1269:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1270:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        1271:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h7A;
        end
        1272:
        begin
            RED=8'hC0;
            GRN=8'hA9;
            BLU=8'h7C;
        end
        1273:
        begin
            RED=8'h81;
            GRN=8'h80;
            BLU=8'h5C;
        end
        1274:
        begin
            RED=8'h4D;
            GRN=8'h50;
            BLU=8'h3E;
        end
        1275:
        begin
            RED=8'h2F;
            GRN=8'h31;
            BLU=8'h2A;
        end
        1276:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1277:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1278:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1279:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1280:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1281:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1282:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1283:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1284:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1285:
        begin
            RED=8'h80;
            GRN=8'h82;
            BLU=8'h63;
        end
        1286:
        begin
            RED=8'h7E;
            GRN=8'h84;
            BLU=8'h64;
        end
        1287:
        begin
            RED=8'h7B;
            GRN=8'h83;
            BLU=8'h68;
        end
        1288:
        begin
            RED=8'h6E;
            GRN=8'h78;
            BLU=8'h60;
        end
        1289:
        begin
            RED=8'h65;
            GRN=8'h75;
            BLU=8'h5D;
        end
        1290:
        begin
            RED=8'h66;
            GRN=8'h6D;
            BLU=8'h55;
        end
        1291:
        begin
            RED=8'h98;
            GRN=8'h90;
            BLU=8'h73;
        end
        1292:
        begin
            RED=8'hAC;
            GRN=8'h9E;
            BLU=8'h78;
        end
        1293:
        begin
            RED=8'hBE;
            GRN=8'hAF;
            BLU=8'h81;
        end
        1294:
        begin
            RED=8'hD3;
            GRN=8'hB7;
            BLU=8'h84;
        end
        1295:
        begin
            RED=8'hE2;
            GRN=8'hC1;
            BLU=8'h8B;
        end
        1296:
        begin
            RED=8'hE9;
            GRN=8'hC2;
            BLU=8'h88;
        end
        1297:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h84;
        end
        1298:
        begin
            RED=8'hEE;
            GRN=8'hC3;
            BLU=8'h80;
        end
        1299:
        begin
            RED=8'hD2;
            GRN=8'hAB;
            BLU=8'h69;
        end
        1300:
        begin
            RED=8'hE6;
            GRN=8'hC1;
            BLU=8'h85;
        end
        1301:
        begin
            RED=8'hE4;
            GRN=8'hBD;
            BLU=8'h82;
        end
        1302:
        begin
            RED=8'hDC;
            GRN=8'hB2;
            BLU=8'h74;
        end
        1303:
        begin
            RED=8'hCA;
            GRN=8'hB6;
            BLU=8'h7D;
        end
        1304:
        begin
            RED=8'hB7;
            GRN=8'hB4;
            BLU=8'h97;
        end
        1305:
        begin
            RED=8'hBB;
            GRN=8'hCD;
            BLU=8'hC6;
        end
        1306:
        begin
            RED=8'hB8;
            GRN=8'hD9;
            BLU=8'hD2;
        end
        1307:
        begin
            RED=8'hB6;
            GRN=8'hDA;
            BLU=8'hD4;
        end
        1308:
        begin
            RED=8'hBA;
            GRN=8'hD7;
            BLU=8'hD6;
        end
        1309:
        begin
            RED=8'hB7;
            GRN=8'hCC;
            BLU=8'hC0;
        end
        1310:
        begin
            RED=8'h99;
            GRN=8'hA3;
            BLU=8'h8C;
        end
        1311:
        begin
            RED=8'h8F;
            GRN=8'h8F;
            BLU=8'h70;
        end
        1312:
        begin
            RED=8'hAE;
            GRN=8'hA5;
            BLU=8'h79;
        end
        1313:
        begin
            RED=8'hD3;
            GRN=8'hB9;
            BLU=8'h8A;
        end
        1314:
        begin
            RED=8'hE7;
            GRN=8'hBC;
            BLU=8'h8A;
        end
        1315:
        begin
            RED=8'hDC;
            GRN=8'hAD;
            BLU=8'h76;
        end
        1316:
        begin
            RED=8'hD0;
            GRN=8'hA4;
            BLU=8'h6B;
        end
        1317:
        begin
            RED=8'hD4;
            GRN=8'hAC;
            BLU=8'h6F;
        end
        1318:
        begin
            RED=8'hD3;
            GRN=8'hAB;
            BLU=8'h67;
        end
        1319:
        begin
            RED=8'hE6;
            GRN=8'hBD;
            BLU=8'h78;
        end
        1320:
        begin
            RED=8'hF0;
            GRN=8'hC2;
            BLU=8'h84;
        end
        1321:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        1322:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1323:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1324:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1325:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1326:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1327:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1328:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1329:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1330:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1331:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1332:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1333:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1334:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        1335:
        begin
            RED=8'hE4;
            GRN=8'hC1;
            BLU=8'h84;
        end
        1336:
        begin
            RED=8'h95;
            GRN=8'h86;
            BLU=8'h5F;
        end
        1337:
        begin
            RED=8'h80;
            GRN=8'h82;
            BLU=8'h61;
        end
        1338:
        begin
            RED=8'h4E;
            GRN=8'h52;
            BLU=8'h40;
        end
        1339:
        begin
            RED=8'h31;
            GRN=8'h32;
            BLU=8'h2C;
        end
        1340:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1341:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1342:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1343:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1344:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1345:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1346:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1347:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1348:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1349:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h68;
        end
        1350:
        begin
            RED=8'h71;
            GRN=8'h7C;
            BLU=8'h68;
        end
        1351:
        begin
            RED=8'h7E;
            GRN=8'h8E;
            BLU=8'h80;
        end
        1352:
        begin
            RED=8'hA9;
            GRN=8'hBE;
            BLU=8'hAF;
        end
        1353:
        begin
            RED=8'hB1;
            GRN=8'hCE;
            BLU=8'hC5;
        end
        1354:
        begin
            RED=8'hB5;
            GRN=8'hD2;
            BLU=8'hCC;
        end
        1355:
        begin
            RED=8'hB0;
            GRN=8'hCA;
            BLU=8'hC2;
        end
        1356:
        begin
            RED=8'h95;
            GRN=8'hAD;
            BLU=8'hA2;
        end
        1357:
        begin
            RED=8'h91;
            GRN=8'hA9;
            BLU=8'h9D;
        end
        1358:
        begin
            RED=8'h9B;
            GRN=8'hB2;
            BLU=8'hA5;
        end
        1359:
        begin
            RED=8'h95;
            GRN=8'hA3;
            BLU=8'h8B;
        end
        1360:
        begin
            RED=8'hA9;
            GRN=8'hA5;
            BLU=8'h7E;
        end
        1361:
        begin
            RED=8'hD0;
            GRN=8'hB7;
            BLU=8'h84;
        end
        1362:
        begin
            RED=8'hE2;
            GRN=8'hC2;
            BLU=8'h8A;
        end
        1363:
        begin
            RED=8'hC9;
            GRN=8'hA3;
            BLU=8'h67;
        end
        1364:
        begin
            RED=8'hE8;
            GRN=8'hBE;
            BLU=8'h7F;
        end
        1365:
        begin
            RED=8'hDF;
            GRN=8'hBE;
            BLU=8'h87;
        end
        1366:
        begin
            RED=8'hB6;
            GRN=8'hA8;
            BLU=8'h7D;
        end
        1367:
        begin
            RED=8'hA9;
            GRN=8'hC0;
            BLU=8'hAF;
        end
        1368:
        begin
            RED=8'hB9;
            GRN=8'hD8;
            BLU=8'hD4;
        end
        1369:
        begin
            RED=8'hB5;
            GRN=8'hD8;
            BLU=8'hD8;
        end
        1370:
        begin
            RED=8'hB7;
            GRN=8'hDA;
            BLU=8'hCF;
        end
        1371:
        begin
            RED=8'hB9;
            GRN=8'hD9;
            BLU=8'hCD;
        end
        1372:
        begin
            RED=8'hB9;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1373:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hD4;
        end
        1374:
        begin
            RED=8'hB6;
            GRN=8'hDD;
            BLU=8'hD8;
        end
        1375:
        begin
            RED=8'hAA;
            GRN=8'hD4;
            BLU=8'hCF;
        end
        1376:
        begin
            RED=8'h84;
            GRN=8'hA6;
            BLU=8'h9E;
        end
        1377:
        begin
            RED=8'h93;
            GRN=8'hA8;
            BLU=8'h9A;
        end
        1378:
        begin
            RED=8'h8C;
            GRN=8'h8B;
            BLU=8'h6E;
        end
        1379:
        begin
            RED=8'hCA;
            GRN=8'hB1;
            BLU=8'h83;
        end
        1380:
        begin
            RED=8'hE3;
            GRN=8'hBF;
            BLU=8'h89;
        end
        1381:
        begin
            RED=8'hE6;
            GRN=8'hC2;
            BLU=8'h89;
        end
        1382:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h82;
        end
        1383:
        begin
            RED=8'hED;
            GRN=8'hBE;
            BLU=8'h7C;
        end
        1384:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h80;
        end
        1385:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1386:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1387:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1388:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1389:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1390:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1391:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1392:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1393:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1394:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1395:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1396:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1397:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1398:
        begin
            RED=8'hEB;
            GRN=8'hC1;
            BLU=8'h81;
        end
        1399:
        begin
            RED=8'hCF;
            GRN=8'hB7;
            BLU=8'h84;
        end
        1400:
        begin
            RED=8'h82;
            GRN=8'h7B;
            BLU=8'h5C;
        end
        1401:
        begin
            RED=8'h7C;
            GRN=8'h83;
            BLU=8'h65;
        end
        1402:
        begin
            RED=8'h4F;
            GRN=8'h54;
            BLU=8'h43;
        end
        1403:
        begin
            RED=8'h30;
            GRN=8'h30;
            BLU=8'h2A;
        end
        1404:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1405:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1406:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1407:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1408:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1409:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1410:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1411:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1412:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h66;
        end
        1413:
        begin
            RED=8'h71;
            GRN=8'h80;
            BLU=8'h6A;
        end
        1414:
        begin
            RED=8'hA9;
            GRN=8'hBB;
            BLU=8'hB1;
        end
        1415:
        begin
            RED=8'hBB;
            GRN=8'hD4;
            BLU=8'hCF;
        end
        1416:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD1;
        end
        1417:
        begin
            RED=8'hB9;
            GRN=8'hD8;
            BLU=8'hD2;
        end
        1418:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD2;
        end
        1419:
        begin
            RED=8'hB5;
            GRN=8'hD7;
            BLU=8'hD3;
        end
        1420:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hD5;
        end
        1421:
        begin
            RED=8'hA5;
            GRN=8'hC8;
            BLU=8'hC7;
        end
        1422:
        begin
            RED=8'h81;
            GRN=8'hAA;
            BLU=8'hA7;
        end
        1423:
        begin
            RED=8'h94;
            GRN=8'hC1;
            BLU=8'hB7;
        end
        1424:
        begin
            RED=8'h99;
            GRN=8'hC2;
            BLU=8'hB3;
        end
        1425:
        begin
            RED=8'h96;
            GRN=8'hB2;
            BLU=8'hA2;
        end
        1426:
        begin
            RED=8'h98;
            GRN=8'h97;
            BLU=8'h7A;
        end
        1427:
        begin
            RED=8'hD7;
            GRN=8'hB3;
            BLU=8'h7A;
        end
        1428:
        begin
            RED=8'hF3;
            GRN=8'hBE;
            BLU=8'h78;
        end
        1429:
        begin
            RED=8'hD8;
            GRN=8'hBF;
            BLU=8'h8C;
        end
        1430:
        begin
            RED=8'hA2;
            GRN=8'hB3;
            BLU=8'hA0;
        end
        1431:
        begin
            RED=8'hBB;
            GRN=8'hD8;
            BLU=8'hD5;
        end
        1432:
        begin
            RED=8'hB7;
            GRN=8'hDA;
            BLU=8'hD2;
        end
        1433:
        begin
            RED=8'hB3;
            GRN=8'hDC;
            BLU=8'hCE;
        end
        1434:
        begin
            RED=8'hB5;
            GRN=8'hDA;
            BLU=8'hD0;
        end
        1435:
        begin
            RED=8'hB5;
            GRN=8'hD9;
            BLU=8'hD4;
        end
        1436:
        begin
            RED=8'hB5;
            GRN=8'hD9;
            BLU=8'hD4;
        end
        1437:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hD2;
        end
        1438:
        begin
            RED=8'hB9;
            GRN=8'hDA;
            BLU=8'hD0;
        end
        1439:
        begin
            RED=8'hB8;
            GRN=8'hDA;
            BLU=8'hCD;
        end
        1440:
        begin
            RED=8'hB7;
            GRN=8'hD2;
            BLU=8'hD1;
        end
        1441:
        begin
            RED=8'h8A;
            GRN=8'hB5;
            BLU=8'hB1;
        end
        1442:
        begin
            RED=8'h8F;
            GRN=8'hC0;
            BLU=8'hB5;
        end
        1443:
        begin
            RED=8'h94;
            GRN=8'hB1;
            BLU=8'h9E;
        end
        1444:
        begin
            RED=8'h9A;
            GRN=8'h9A;
            BLU=8'h7C;
        end
        1445:
        begin
            RED=8'hD2;
            GRN=8'hB5;
            BLU=8'h83;
        end
        1446:
        begin
            RED=8'hEB;
            GRN=8'hC1;
            BLU=8'h86;
        end
        1447:
        begin
            RED=8'hF3;
            GRN=8'hC0;
            BLU=8'h80;
        end
        1448:
        begin
            RED=8'hEC;
            GRN=8'hBE;
            BLU=8'h7D;
        end
        1449:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1450:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1451:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1452:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1453:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1454:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1455:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1456:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1457:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1458:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1459:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        1460:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        1461:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1462:
        begin
            RED=8'hE9;
            GRN=8'hC1;
            BLU=8'h83;
        end
        1463:
        begin
            RED=8'h9C;
            GRN=8'h8D;
            BLU=8'h61;
        end
        1464:
        begin
            RED=8'h7E;
            GRN=8'h7D;
            BLU=8'h62;
        end
        1465:
        begin
            RED=8'h7B;
            GRN=8'h84;
            BLU=8'h68;
        end
        1466:
        begin
            RED=8'h4F;
            GRN=8'h53;
            BLU=8'h43;
        end
        1467:
        begin
            RED=8'h30;
            GRN=8'h30;
            BLU=8'h29;
        end
        1468:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1469:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1470:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1471:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1472:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h62;
        end
        1473:
        begin
            RED=8'h80;
            GRN=8'h82;
            BLU=8'h64;
        end
        1474:
        begin
            RED=8'h83;
            GRN=8'h82;
            BLU=8'h68;
        end
        1475:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h67;
        end
        1476:
        begin
            RED=8'h74;
            GRN=8'h81;
            BLU=8'h66;
        end
        1477:
        begin
            RED=8'h98;
            GRN=8'hB4;
            BLU=8'hAB;
        end
        1478:
        begin
            RED=8'hBA;
            GRN=8'hD8;
            BLU=8'hCF;
        end
        1479:
        begin
            RED=8'hB7;
            GRN=8'hDA;
            BLU=8'hD1;
        end
        1480:
        begin
            RED=8'hB1;
            GRN=8'hD8;
            BLU=8'hCD;
        end
        1481:
        begin
            RED=8'hB5;
            GRN=8'hD8;
            BLU=8'hD1;
        end
        1482:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1483:
        begin
            RED=8'hB9;
            GRN=8'hD9;
            BLU=8'hD4;
        end
        1484:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1485:
        begin
            RED=8'hB7;
            GRN=8'hD9;
            BLU=8'hD4;
        end
        1486:
        begin
            RED=8'h9F;
            GRN=8'hC9;
            BLU=8'hC3;
        end
        1487:
        begin
            RED=8'h87;
            GRN=8'hB2;
            BLU=8'hAB;
        end
        1488:
        begin
            RED=8'h93;
            GRN=8'hC0;
            BLU=8'hB9;
        end
        1489:
        begin
            RED=8'h93;
            GRN=8'hC0;
            BLU=8'hB9;
        end
        1490:
        begin
            RED=8'h96;
            GRN=8'hB2;
            BLU=8'hA5;
        end
        1491:
        begin
            RED=8'hD3;
            GRN=8'hB7;
            BLU=8'h86;
        end
        1492:
        begin
            RED=8'hF3;
            GRN=8'hBD;
            BLU=8'h7A;
        end
        1493:
        begin
            RED=8'hB2;
            GRN=8'hAC;
            BLU=8'h88;
        end
        1494:
        begin
            RED=8'hB6;
            GRN=8'hD7;
            BLU=8'hCC;
        end
        1495:
        begin
            RED=8'hB7;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1496:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD2;
        end
        1497:
        begin
            RED=8'hB8;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        1498:
        begin
            RED=8'hA8;
            GRN=8'hC9;
            BLU=8'hC4;
        end
        1499:
        begin
            RED=8'hAD;
            GRN=8'hCD;
            BLU=8'hC9;
        end
        1500:
        begin
            RED=8'hB8;
            GRN=8'hD9;
            BLU=8'hD4;
        end
        1501:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD2;
        end
        1502:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1503:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD2;
        end
        1504:
        begin
            RED=8'hB6;
            GRN=8'hD8;
            BLU=8'hD2;
        end
        1505:
        begin
            RED=8'hAB;
            GRN=8'hCD;
            BLU=8'hC8;
        end
        1506:
        begin
            RED=8'h8B;
            GRN=8'hB3;
            BLU=8'hAC;
        end
        1507:
        begin
            RED=8'h91;
            GRN=8'hC1;
            BLU=8'hB7;
        end
        1508:
        begin
            RED=8'h92;
            GRN=8'hC0;
            BLU=8'hB3;
        end
        1509:
        begin
            RED=8'h98;
            GRN=8'hAC;
            BLU=8'h9A;
        end
        1510:
        begin
            RED=8'hBA;
            GRN=8'hA8;
            BLU=8'h81;
        end
        1511:
        begin
            RED=8'hF1;
            GRN=8'hBE;
            BLU=8'h7D;
        end
        1512:
        begin
            RED=8'hEC;
            GRN=8'hC1;
            BLU=8'h7B;
        end
        1513:
        begin
            RED=8'hEB;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1514:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1515:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1516:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1517:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1518:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1519:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1520:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1521:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1522:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h81;
        end
        1523:
        begin
            RED=8'hF0;
            GRN=8'hBF;
            BLU=8'h7C;
        end
        1524:
        begin
            RED=8'hF2;
            GRN=8'hBF;
            BLU=8'h78;
        end
        1525:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h81;
        end
        1526:
        begin
            RED=8'hD7;
            GRN=8'hBB;
            BLU=8'h87;
        end
        1527:
        begin
            RED=8'h79;
            GRN=8'h7B;
            BLU=8'h5A;
        end
        1528:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h63;
        end
        1529:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h69;
        end
        1530:
        begin
            RED=8'h50;
            GRN=8'h53;
            BLU=8'h44;
        end
        1531:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h28;
        end
        1532:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1533:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1534:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1535:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1536:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h64;
        end
        1537:
        begin
            RED=8'h80;
            GRN=8'h82;
            BLU=8'h63;
        end
        1538:
        begin
            RED=8'h81;
            GRN=8'h82;
            BLU=8'h66;
        end
        1539:
        begin
            RED=8'h7C;
            GRN=8'h82;
            BLU=8'h67;
        end
        1540:
        begin
            RED=8'h77;
            GRN=8'h87;
            BLU=8'h70;
        end
        1541:
        begin
            RED=8'hB8;
            GRN=8'hD7;
            BLU=8'hCE;
        end
        1542:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD0;
        end
        1543:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hD0;
        end
        1544:
        begin
            RED=8'hA6;
            GRN=8'hCB;
            BLU=8'hC0;
        end
        1545:
        begin
            RED=8'hA5;
            GRN=8'hC7;
            BLU=8'hC0;
        end
        1546:
        begin
            RED=8'hB7;
            GRN=8'hD7;
            BLU=8'hD2;
        end
        1547:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1548:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1549:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1550:
        begin
            RED=8'hB9;
            GRN=8'hDA;
            BLU=8'hD5;
        end
        1551:
        begin
            RED=8'h8D;
            GRN=8'hB3;
            BLU=8'hAC;
        end
        1552:
        begin
            RED=8'h92;
            GRN=8'hC0;
            BLU=8'hB6;
        end
        1553:
        begin
            RED=8'h90;
            GRN=8'hC2;
            BLU=8'hB7;
        end
        1554:
        begin
            RED=8'h93;
            GRN=8'hBF;
            BLU=8'hB6;
        end
        1555:
        begin
            RED=8'hA9;
            GRN=8'hA1;
            BLU=8'h7B;
        end
        1556:
        begin
            RED=8'hE5;
            GRN=8'hC1;
            BLU=8'h8B;
        end
        1557:
        begin
            RED=8'hAD;
            GRN=8'hAF;
            BLU=8'h99;
        end
        1558:
        begin
            RED=8'hBA;
            GRN=8'hD9;
            BLU=8'hD2;
        end
        1559:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1560:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1561:
        begin
            RED=8'hB7;
            GRN=8'hD7;
            BLU=8'hD2;
        end
        1562:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1563:
        begin
            RED=8'h9D;
            GRN=8'hBD;
            BLU=8'hB8;
        end
        1564:
        begin
            RED=8'hB0;
            GRN=8'hD0;
            BLU=8'hCB;
        end
        1565:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1566:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1567:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1568:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        1569:
        begin
            RED=8'hB6;
            GRN=8'hD7;
            BLU=8'hD2;
        end
        1570:
        begin
            RED=8'h89;
            GRN=8'hAF;
            BLU=8'hA8;
        end
        1571:
        begin
            RED=8'h90;
            GRN=8'hC0;
            BLU=8'hB6;
        end
        1572:
        begin
            RED=8'h8C;
            GRN=8'hC1;
            BLU=8'hB8;
        end
        1573:
        begin
            RED=8'h95;
            GRN=8'hC0;
            BLU=8'hBB;
        end
        1574:
        begin
            RED=8'h97;
            GRN=8'h9D;
            BLU=8'h83;
        end
        1575:
        begin
            RED=8'hE5;
            GRN=8'hC0;
            BLU=8'h85;
        end
        1576:
        begin
            RED=8'hEF;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        1577:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1578:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1579:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1580:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1581:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1582:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1583:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1584:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1585:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1586:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h81;
        end
        1587:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h7C;
        end
        1588:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h7B;
        end
        1589:
        begin
            RED=8'hE6;
            GRN=8'hC2;
            BLU=8'h87;
        end
        1590:
        begin
            RED=8'hA6;
            GRN=8'h91;
            BLU=8'h63;
        end
        1591:
        begin
            RED=8'h7C;
            GRN=8'h80;
            BLU=8'h61;
        end
        1592:
        begin
            RED=8'h7D;
            GRN=8'h82;
            BLU=8'h62;
        end
        1593:
        begin
            RED=8'h7D;
            GRN=8'h81;
            BLU=8'h68;
        end
        1594:
        begin
            RED=8'h50;
            GRN=8'h53;
            BLU=8'h44;
        end
        1595:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h28;
        end
        1596:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1597:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1598:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1599:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1600:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h66;
        end
        1601:
        begin
            RED=8'h80;
            GRN=8'h82;
            BLU=8'h63;
        end
        1602:
        begin
            RED=8'h7F;
            GRN=8'h82;
            BLU=8'h63;
        end
        1603:
        begin
            RED=8'h7A;
            GRN=8'h85;
            BLU=8'h6C;
        end
        1604:
        begin
            RED=8'h9E;
            GRN=8'hB3;
            BLU=8'hA3;
        end
        1605:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hCF;
        end
        1606:
        begin
            RED=8'hB7;
            GRN=8'hDA;
            BLU=8'hD0;
        end
        1607:
        begin
            RED=8'hB8;
            GRN=8'hD9;
            BLU=8'hD0;
        end
        1608:
        begin
            RED=8'hB9;
            GRN=8'hDB;
            BLU=8'hD2;
        end
        1609:
        begin
            RED=8'hA2;
            GRN=8'hC3;
            BLU=8'hBD;
        end
        1610:
        begin
            RED=8'hA6;
            GRN=8'hC6;
            BLU=8'hC1;
        end
        1611:
        begin
            RED=8'hB9;
            GRN=8'hD9;
            BLU=8'hD4;
        end
        1612:
        begin
            RED=8'hBA;
            GRN=8'hDA;
            BLU=8'hD5;
        end
        1613:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1614:
        begin
            RED=8'hB9;
            GRN=8'hD6;
            BLU=8'hD1;
        end
        1615:
        begin
            RED=8'hA5;
            GRN=8'hC8;
            BLU=8'hC1;
        end
        1616:
        begin
            RED=8'h90;
            GRN=8'hBC;
            BLU=8'hB2;
        end
        1617:
        begin
            RED=8'h8F;
            GRN=8'hC3;
            BLU=8'hB6;
        end
        1618:
        begin
            RED=8'h92;
            GRN=8'hC0;
            BLU=8'hB4;
        end
        1619:
        begin
            RED=8'h9B;
            GRN=8'h9D;
            BLU=8'h7A;
        end
        1620:
        begin
            RED=8'hCF;
            GRN=8'hBA;
            BLU=8'h90;
        end
        1621:
        begin
            RED=8'hB9;
            GRN=8'hC6;
            BLU=8'hB9;
        end
        1622:
        begin
            RED=8'hB8;
            GRN=8'hD6;
            BLU=8'hD2;
        end
        1623:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1624:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1625:
        begin
            RED=8'hB7;
            GRN=8'hD7;
            BLU=8'hD2;
        end
        1626:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1627:
        begin
            RED=8'hB7;
            GRN=8'hD7;
            BLU=8'hD2;
        end
        1628:
        begin
            RED=8'h9D;
            GRN=8'hBD;
            BLU=8'hB8;
        end
        1629:
        begin
            RED=8'hB2;
            GRN=8'hD2;
            BLU=8'hCD;
        end
        1630:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1631:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1632:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        1633:
        begin
            RED=8'hB7;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1634:
        begin
            RED=8'h96;
            GRN=8'hBC;
            BLU=8'hB5;
        end
        1635:
        begin
            RED=8'h8F;
            GRN=8'hC0;
            BLU=8'hB5;
        end
        1636:
        begin
            RED=8'h8D;
            GRN=8'hC4;
            BLU=8'hBC;
        end
        1637:
        begin
            RED=8'h8C;
            GRN=8'hC4;
            BLU=8'hC4;
        end
        1638:
        begin
            RED=8'h97;
            GRN=8'hB6;
            BLU=8'hA6;
        end
        1639:
        begin
            RED=8'hC7;
            GRN=8'hB4;
            BLU=8'h82;
        end
        1640:
        begin
            RED=8'hEF;
            GRN=8'hC1;
            BLU=8'h80;
        end
        1641:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        1642:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1643:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1644:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1645:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1646:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1647:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1648:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1649:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1650:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h80;
        end
        1651:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        1652:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h80;
        end
        1653:
        begin
            RED=8'hD3;
            GRN=8'hB9;
            BLU=8'h85;
        end
        1654:
        begin
            RED=8'h87;
            GRN=8'h7E;
            BLU=8'h59;
        end
        1655:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h64;
        end
        1656:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1657:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h69;
        end
        1658:
        begin
            RED=8'h52;
            GRN=8'h54;
            BLU=8'h46;
        end
        1659:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1660:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1661:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1662:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1663:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1664:
        begin
            RED=8'h7F;
            GRN=8'h81;
            BLU=8'h68;
        end
        1665:
        begin
            RED=8'h81;
            GRN=8'h82;
            BLU=8'h63;
        end
        1666:
        begin
            RED=8'h7E;
            GRN=8'h85;
            BLU=8'h62;
        end
        1667:
        begin
            RED=8'h73;
            GRN=8'h82;
            BLU=8'h6B;
        end
        1668:
        begin
            RED=8'hA7;
            GRN=8'hC0;
            BLU=8'hB5;
        end
        1669:
        begin
            RED=8'hB5;
            GRN=8'hDB;
            BLU=8'hD0;
        end
        1670:
        begin
            RED=8'hB6;
            GRN=8'hDA;
            BLU=8'hD0;
        end
        1671:
        begin
            RED=8'hB3;
            GRN=8'hD4;
            BLU=8'hCB;
        end
        1672:
        begin
            RED=8'hBA;
            GRN=8'hD8;
            BLU=8'hD0;
        end
        1673:
        begin
            RED=8'hBA;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        1674:
        begin
            RED=8'h9D;
            GRN=8'hBD;
            BLU=8'hB8;
        end
        1675:
        begin
            RED=8'hB1;
            GRN=8'hD1;
            BLU=8'hCC;
        end
        1676:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1677:
        begin
            RED=8'hB7;
            GRN=8'hD8;
            BLU=8'hD2;
        end
        1678:
        begin
            RED=8'hB8;
            GRN=8'hD9;
            BLU=8'hD1;
        end
        1679:
        begin
            RED=8'hAC;
            GRN=8'hD0;
            BLU=8'hC7;
        end
        1680:
        begin
            RED=8'h8D;
            GRN=8'hB6;
            BLU=8'hAB;
        end
        1681:
        begin
            RED=8'h93;
            GRN=8'hC0;
            BLU=8'hB4;
        end
        1682:
        begin
            RED=8'h9C;
            GRN=8'hB7;
            BLU=8'hA4;
        end
        1683:
        begin
            RED=8'h96;
            GRN=8'h86;
            BLU=8'h5C;
        end
        1684:
        begin
            RED=8'hAB;
            GRN=8'h96;
            BLU=8'h6D;
        end
        1685:
        begin
            RED=8'hBB;
            GRN=8'hCF;
            BLU=8'hC5;
        end
        1686:
        begin
            RED=8'hB4;
            GRN=8'hD7;
            BLU=8'hD2;
        end
        1687:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1688:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1689:
        begin
            RED=8'h9C;
            GRN=8'hBC;
            BLU=8'hB7;
        end
        1690:
        begin
            RED=8'hB0;
            GRN=8'hD0;
            BLU=8'hCB;
        end
        1691:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1692:
        begin
            RED=8'hB6;
            GRN=8'hD6;
            BLU=8'hD1;
        end
        1693:
        begin
            RED=8'h9F;
            GRN=8'hBF;
            BLU=8'hBA;
        end
        1694:
        begin
            RED=8'hB3;
            GRN=8'hD3;
            BLU=8'hCE;
        end
        1695:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1696:
        begin
            RED=8'hB7;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        1697:
        begin
            RED=8'hB7;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1698:
        begin
            RED=8'h97;
            GRN=8'hBE;
            BLU=8'hB6;
        end
        1699:
        begin
            RED=8'h8F;
            GRN=8'hC0;
            BLU=8'hB5;
        end
        1700:
        begin
            RED=8'h8E;
            GRN=8'hC3;
            BLU=8'hB7;
        end
        1701:
        begin
            RED=8'h8D;
            GRN=8'hC4;
            BLU=8'hC0;
        end
        1702:
        begin
            RED=8'h94;
            GRN=8'hC1;
            BLU=8'hB4;
        end
        1703:
        begin
            RED=8'hAC;
            GRN=8'hA7;
            BLU=8'h7D;
        end
        1704:
        begin
            RED=8'hEE;
            GRN=8'hC1;
            BLU=8'h85;
        end
        1705:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h7F;
        end
        1706:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1707:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1708:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1709:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1710:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1711:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1712:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1713:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1714:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1715:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        1716:
        begin
            RED=8'hE7;
            GRN=8'hC1;
            BLU=8'h85;
        end
        1717:
        begin
            RED=8'h9D;
            GRN=8'h8C;
            BLU=8'h60;
        end
        1718:
        begin
            RED=8'h80;
            GRN=8'h80;
            BLU=8'h62;
        end
        1719:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        1720:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1721:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h69;
        end
        1722:
        begin
            RED=8'h53;
            GRN=8'h55;
            BLU=8'h47;
        end
        1723:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1724:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1725:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1726:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1727:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1728:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h66;
        end
        1729:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h61;
        end
        1730:
        begin
            RED=8'h7C;
            GRN=8'h83;
            BLU=8'h62;
        end
        1731:
        begin
            RED=8'h70;
            GRN=8'h80;
            BLU=8'h6B;
        end
        1732:
        begin
            RED=8'hA7;
            GRN=8'hC2;
            BLU=8'hB7;
        end
        1733:
        begin
            RED=8'hB4;
            GRN=8'hDA;
            BLU=8'hD2;
        end
        1734:
        begin
            RED=8'hB7;
            GRN=8'hD9;
            BLU=8'hD2;
        end
        1735:
        begin
            RED=8'h9E;
            GRN=8'hBD;
            BLU=8'hB7;
        end
        1736:
        begin
            RED=8'hB3;
            GRN=8'hD3;
            BLU=8'hCB;
        end
        1737:
        begin
            RED=8'hB8;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        1738:
        begin
            RED=8'hB6;
            GRN=8'hD7;
            BLU=8'hD1;
        end
        1739:
        begin
            RED=8'h98;
            GRN=8'hB8;
            BLU=8'hB0;
        end
        1740:
        begin
            RED=8'hB3;
            GRN=8'hD4;
            BLU=8'hCB;
        end
        1741:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hD1;
        end
        1742:
        begin
            RED=8'hB3;
            GRN=8'hDA;
            BLU=8'hD0;
        end
        1743:
        begin
            RED=8'hAC;
            GRN=8'hD3;
            BLU=8'hCC;
        end
        1744:
        begin
            RED=8'h92;
            GRN=8'hAF;
            BLU=8'hA3;
        end
        1745:
        begin
            RED=8'h9C;
            GRN=8'hAA;
            BLU=8'h91;
        end
        1746:
        begin
            RED=8'hB9;
            GRN=8'hB1;
            BLU=8'h89;
        end
        1747:
        begin
            RED=8'hE7;
            GRN=8'hBF;
            BLU=8'h84;
        end
        1748:
        begin
            RED=8'hCC;
            GRN=8'hAD;
            BLU=8'h7E;
        end
        1749:
        begin
            RED=8'hBD;
            GRN=8'hD0;
            BLU=8'hC3;
        end
        1750:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hD0;
        end
        1751:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1752:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1753:
        begin
            RED=8'hB7;
            GRN=8'hD7;
            BLU=8'hD2;
        end
        1754:
        begin
            RED=8'h97;
            GRN=8'hB7;
            BLU=8'hB2;
        end
        1755:
        begin
            RED=8'hAF;
            GRN=8'hCF;
            BLU=8'hCA;
        end
        1756:
        begin
            RED=8'hB9;
            GRN=8'hDB;
            BLU=8'hD5;
        end
        1757:
        begin
            RED=8'hB7;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1758:
        begin
            RED=8'hA0;
            GRN=8'hC2;
            BLU=8'hBC;
        end
        1759:
        begin
            RED=8'hB4;
            GRN=8'hD6;
            BLU=8'hD0;
        end
        1760:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        1761:
        begin
            RED=8'hB9;
            GRN=8'hD9;
            BLU=8'hD4;
        end
        1762:
        begin
            RED=8'h95;
            GRN=8'hBA;
            BLU=8'hB3;
        end
        1763:
        begin
            RED=8'h90;
            GRN=8'hBF;
            BLU=8'hB7;
        end
        1764:
        begin
            RED=8'h8F;
            GRN=8'hC2;
            BLU=8'hB5;
        end
        1765:
        begin
            RED=8'h90;
            GRN=8'hC4;
            BLU=8'hB9;
        end
        1766:
        begin
            RED=8'h93;
            GRN=8'hC2;
            BLU=8'hB6;
        end
        1767:
        begin
            RED=8'h94;
            GRN=8'h94;
            BLU=8'h6F;
        end
        1768:
        begin
            RED=8'hD9;
            GRN=8'hB2;
            BLU=8'h7C;
        end
        1769:
        begin
            RED=8'hE7;
            GRN=8'hBB;
            BLU=8'h82;
        end
        1770:
        begin
            RED=8'hEB;
            GRN=8'hBF;
            BLU=8'h85;
        end
        1771:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h85;
        end
        1772:
        begin
            RED=8'hEB;
            GRN=8'hC0;
            BLU=8'h82;
        end
        1773:
        begin
            RED=8'hEB;
            GRN=8'hC0;
            BLU=8'h81;
        end
        1774:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1775:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h80;
        end
        1776:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h80;
        end
        1777:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1778:
        begin
            RED=8'hF1;
            GRN=8'hC0;
            BLU=8'h7C;
        end
        1779:
        begin
            RED=8'hEC;
            GRN=8'hC1;
            BLU=8'h81;
        end
        1780:
        begin
            RED=8'hCB;
            GRN=8'hB1;
            BLU=8'h7E;
        end
        1781:
        begin
            RED=8'h81;
            GRN=8'h7B;
            BLU=8'h56;
        end
        1782:
        begin
            RED=8'h7C;
            GRN=8'h82;
            BLU=8'h66;
        end
        1783:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        1784:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1785:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h69;
        end
        1786:
        begin
            RED=8'h54;
            GRN=8'h56;
            BLU=8'h48;
        end
        1787:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h28;
        end
        1788:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1789:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1790:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1791:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1792:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h62;
        end
        1793:
        begin
            RED=8'h7E;
            GRN=8'h84;
            BLU=8'h60;
        end
        1794:
        begin
            RED=8'h7C;
            GRN=8'h82;
            BLU=8'h63;
        end
        1795:
        begin
            RED=8'h76;
            GRN=8'h83;
            BLU=8'h6C;
        end
        1796:
        begin
            RED=8'hA0;
            GRN=8'hB6;
            BLU=8'hA9;
        end
        1797:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        1798:
        begin
            RED=8'hB7;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1799:
        begin
            RED=8'hB7;
            GRN=8'hD7;
            BLU=8'hD2;
        end
        1800:
        begin
            RED=8'h93;
            GRN=8'hB4;
            BLU=8'hAD;
        end
        1801:
        begin
            RED=8'hB3;
            GRN=8'hD6;
            BLU=8'hCF;
        end
        1802:
        begin
            RED=8'hBB;
            GRN=8'hDD;
            BLU=8'hD6;
        end
        1803:
        begin
            RED=8'hB6;
            GRN=8'hD7;
            BLU=8'hD0;
        end
        1804:
        begin
            RED=8'hAA;
            GRN=8'hCE;
            BLU=8'hC5;
        end
        1805:
        begin
            RED=8'hB5;
            GRN=8'hDB;
            BLU=8'hD1;
        end
        1806:
        begin
            RED=8'hB6;
            GRN=8'hDA;
            BLU=8'hCE;
        end
        1807:
        begin
            RED=8'hAF;
            GRN=8'hC5;
            BLU=8'hB7;
        end
        1808:
        begin
            RED=8'h93;
            GRN=8'h92;
            BLU=8'h76;
        end
        1809:
        begin
            RED=8'hDA;
            GRN=8'hC0;
            BLU=8'h8D;
        end
        1810:
        begin
            RED=8'hE6;
            GRN=8'hC3;
            BLU=8'h82;
        end
        1811:
        begin
            RED=8'hF1;
            GRN=8'hC0;
            BLU=8'h79;
        end
        1812:
        begin
            RED=8'hDD;
            GRN=8'hBA;
            BLU=8'h85;
        end
        1813:
        begin
            RED=8'hB9;
            GRN=8'hC5;
            BLU=8'hB3;
        end
        1814:
        begin
            RED=8'hB7;
            GRN=8'hD7;
            BLU=8'hCF;
        end
        1815:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1816:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1817:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1818:
        begin
            RED=8'hB4;
            GRN=8'hD4;
            BLU=8'hCF;
        end
        1819:
        begin
            RED=8'h99;
            GRN=8'hBA;
            BLU=8'hB5;
        end
        1820:
        begin
            RED=8'hAF;
            GRN=8'hD2;
            BLU=8'hCC;
        end
        1821:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        1822:
        begin
            RED=8'hB5;
            GRN=8'hD8;
            BLU=8'hD2;
        end
        1823:
        begin
            RED=8'hB5;
            GRN=8'hD8;
            BLU=8'hD2;
        end
        1824:
        begin
            RED=8'hB6;
            GRN=8'hDA;
            BLU=8'hD3;
        end
        1825:
        begin
            RED=8'hB6;
            GRN=8'hD7;
            BLU=8'hD1;
        end
        1826:
        begin
            RED=8'h8A;
            GRN=8'hAE;
            BLU=8'hA9;
        end
        1827:
        begin
            RED=8'h94;
            GRN=8'hC3;
            BLU=8'hBD;
        end
        1828:
        begin
            RED=8'h8E;
            GRN=8'hC4;
            BLU=8'hB8;
        end
        1829:
        begin
            RED=8'h8E;
            GRN=8'hC5;
            BLU=8'hBA;
        end
        1830:
        begin
            RED=8'h96;
            GRN=8'hC0;
            BLU=8'hB4;
        end
        1831:
        begin
            RED=8'hAB;
            GRN=8'hA5;
            BLU=8'h81;
        end
        1832:
        begin
            RED=8'hD8;
            GRN=8'hB2;
            BLU=8'h7E;
        end
        1833:
        begin
            RED=8'hD0;
            GRN=8'hA7;
            BLU=8'h72;
        end
        1834:
        begin
            RED=8'hC0;
            GRN=8'h97;
            BLU=8'h62;
        end
        1835:
        begin
            RED=8'hC3;
            GRN=8'h9A;
            BLU=8'h61;
        end
        1836:
        begin
            RED=8'hD8;
            GRN=8'hB0;
            BLU=8'h74;
        end
        1837:
        begin
            RED=8'hE7;
            GRN=8'hBF;
            BLU=8'h82;
        end
        1838:
        begin
            RED=8'hE9;
            GRN=8'hC0;
            BLU=8'h80;
        end
        1839:
        begin
            RED=8'hEA;
            GRN=8'hC0;
            BLU=8'h81;
        end
        1840:
        begin
            RED=8'hE9;
            GRN=8'hC0;
            BLU=8'h80;
        end
        1841:
        begin
            RED=8'hEC;
            GRN=8'hC2;
            BLU=8'h82;
        end
        1842:
        begin
            RED=8'hEF;
            GRN=8'hBE;
            BLU=8'h78;
        end
        1843:
        begin
            RED=8'hE5;
            GRN=8'hBF;
            BLU=8'h85;
        end
        1844:
        begin
            RED=8'h8F;
            GRN=8'h84;
            BLU=8'h5B;
        end
        1845:
        begin
            RED=8'h7F;
            GRN=8'h84;
            BLU=8'h64;
        end
        1846:
        begin
            RED=8'h7A;
            GRN=8'h82;
            BLU=8'h63;
        end
        1847:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        1848:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1849:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h69;
        end
        1850:
        begin
            RED=8'h55;
            GRN=8'h57;
            BLU=8'h4A;
        end
        1851:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h28;
        end
        1852:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1853:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1854:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1855:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1856:
        begin
            RED=8'h7C;
            GRN=8'h85;
            BLU=8'h63;
        end
        1857:
        begin
            RED=8'h7E;
            GRN=8'h84;
            BLU=8'h61;
        end
        1858:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h61;
        end
        1859:
        begin
            RED=8'h7A;
            GRN=8'h83;
            BLU=8'h6A;
        end
        1860:
        begin
            RED=8'h7B;
            GRN=8'h8D;
            BLU=8'h7B;
        end
        1861:
        begin
            RED=8'hBA;
            GRN=8'hD7;
            BLU=8'hCE;
        end
        1862:
        begin
            RED=8'hB8;
            GRN=8'hD9;
            BLU=8'hD0;
        end
        1863:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hD1;
        end
        1864:
        begin
            RED=8'hB3;
            GRN=8'hD4;
            BLU=8'hCE;
        end
        1865:
        begin
            RED=8'h95;
            GRN=8'hB4;
            BLU=8'hAC;
        end
        1866:
        begin
            RED=8'hB5;
            GRN=8'hD7;
            BLU=8'hD0;
        end
        1867:
        begin
            RED=8'hB4;
            GRN=8'hD9;
            BLU=8'hD6;
        end
        1868:
        begin
            RED=8'hB4;
            GRN=8'hDA;
            BLU=8'hD7;
        end
        1869:
        begin
            RED=8'hB5;
            GRN=8'hD7;
            BLU=8'hD1;
        end
        1870:
        begin
            RED=8'hBA;
            GRN=8'hCA;
            BLU=8'hB3;
        end
        1871:
        begin
            RED=8'hB7;
            GRN=8'hA8;
            BLU=8'h80;
        end
        1872:
        begin
            RED=8'hE6;
            GRN=8'hBF;
            BLU=8'h86;
        end
        1873:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h80;
        end
        1874:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        1875:
        begin
            RED=8'hF0;
            GRN=8'hC0;
            BLU=8'h7C;
        end
        1876:
        begin
            RED=8'hE5;
            GRN=8'hC1;
            BLU=8'h8A;
        end
        1877:
        begin
            RED=8'hAB;
            GRN=8'hAE;
            BLU=8'h92;
        end
        1878:
        begin
            RED=8'hBA;
            GRN=8'hD9;
            BLU=8'hD1;
        end
        1879:
        begin
            RED=8'hB8;
            GRN=8'hD9;
            BLU=8'hD4;
        end
        1880:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1881:
        begin
            RED=8'hB7;
            GRN=8'hD7;
            BLU=8'hD2;
        end
        1882:
        begin
            RED=8'hB9;
            GRN=8'hD9;
            BLU=8'hD4;
        end
        1883:
        begin
            RED=8'hB5;
            GRN=8'hD7;
            BLU=8'hD1;
        end
        1884:
        begin
            RED=8'hA1;
            GRN=8'hC4;
            BLU=8'hBE;
        end
        1885:
        begin
            RED=8'hB4;
            GRN=8'hD7;
            BLU=8'hD1;
        end
        1886:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        1887:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        1888:
        begin
            RED=8'hB9;
            GRN=8'hDB;
            BLU=8'hD4;
        end
        1889:
        begin
            RED=8'hB1;
            GRN=8'hD6;
            BLU=8'hCF;
        end
        1890:
        begin
            RED=8'h80;
            GRN=8'hAA;
            BLU=8'hA3;
        end
        1891:
        begin
            RED=8'h8F;
            GRN=8'hC2;
            BLU=8'hBA;
        end
        1892:
        begin
            RED=8'h8C;
            GRN=8'hC3;
            BLU=8'hBB;
        end
        1893:
        begin
            RED=8'h8D;
            GRN=8'hC4;
            BLU=8'hBE;
        end
        1894:
        begin
            RED=8'h9B;
            GRN=8'hB9;
            BLU=8'hA8;
        end
        1895:
        begin
            RED=8'hC7;
            GRN=8'hB3;
            BLU=8'h84;
        end
        1896:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h82;
        end
        1897:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h85;
        end
        1898:
        begin
            RED=8'hEA;
            GRN=8'hC0;
            BLU=8'h85;
        end
        1899:
        begin
            RED=8'hEB;
            GRN=8'hC1;
            BLU=8'h85;
        end
        1900:
        begin
            RED=8'hE4;
            GRN=8'hBA;
            BLU=8'h7E;
        end
        1901:
        begin
            RED=8'hD4;
            GRN=8'hAA;
            BLU=8'h6E;
        end
        1902:
        begin
            RED=8'hC9;
            GRN=8'hA1;
            BLU=8'h64;
        end
        1903:
        begin
            RED=8'hCC;
            GRN=8'hA4;
            BLU=8'h67;
        end
        1904:
        begin
            RED=8'hDA;
            GRN=8'hB2;
            BLU=8'h75;
        end
        1905:
        begin
            RED=8'hE5;
            GRN=8'hBD;
            BLU=8'h80;
        end
        1906:
        begin
            RED=8'hE8;
            GRN=8'hC2;
            BLU=8'h87;
        end
        1907:
        begin
            RED=8'hB8;
            GRN=8'hA0;
            BLU=8'h6F;
        end
        1908:
        begin
            RED=8'h82;
            GRN=8'h80;
            BLU=8'h5C;
        end
        1909:
        begin
            RED=8'h7F;
            GRN=8'h85;
            BLU=8'h66;
        end
        1910:
        begin
            RED=8'h7F;
            GRN=8'h85;
            BLU=8'h65;
        end
        1911:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        1912:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1913:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h69;
        end
        1914:
        begin
            RED=8'h55;
            GRN=8'h57;
            BLU=8'h4A;
        end
        1915:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h28;
        end
        1916:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1917:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1918:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1919:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1920:
        begin
            RED=8'h7B;
            GRN=8'h85;
            BLU=8'h64;
        end
        1921:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h61;
        end
        1922:
        begin
            RED=8'h81;
            GRN=8'h82;
            BLU=8'h61;
        end
        1923:
        begin
            RED=8'h7D;
            GRN=8'h82;
            BLU=8'h65;
        end
        1924:
        begin
            RED=8'h74;
            GRN=8'h7F;
            BLU=8'h69;
        end
        1925:
        begin
            RED=8'hA9;
            GRN=8'hBD;
            BLU=8'hB1;
        end
        1926:
        begin
            RED=8'hB8;
            GRN=8'hD9;
            BLU=8'hCC;
        end
        1927:
        begin
            RED=8'hB4;
            GRN=8'hDB;
            BLU=8'hD0;
        end
        1928:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1929:
        begin
            RED=8'hB5;
            GRN=8'hD4;
            BLU=8'hCC;
        end
        1930:
        begin
            RED=8'hB4;
            GRN=8'hD8;
            BLU=8'hD1;
        end
        1931:
        begin
            RED=8'hB3;
            GRN=8'hD9;
            BLU=8'hD7;
        end
        1932:
        begin
            RED=8'hBC;
            GRN=8'hD8;
            BLU=8'hD4;
        end
        1933:
        begin
            RED=8'hB8;
            GRN=8'hC5;
            BLU=8'hB7;
        end
        1934:
        begin
            RED=8'hBC;
            GRN=8'hAC;
            BLU=8'h83;
        end
        1935:
        begin
            RED=8'hEA;
            GRN=8'hC0;
            BLU=8'h88;
        end
        1936:
        begin
            RED=8'hF5;
            GRN=8'hBD;
            BLU=8'h78;
        end
        1937:
        begin
            RED=8'hF0;
            GRN=8'hC0;
            BLU=8'h79;
        end
        1938:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        1939:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h80;
        end
        1940:
        begin
            RED=8'hE8;
            GRN=8'hC2;
            BLU=8'h82;
        end
        1941:
        begin
            RED=8'hCD;
            GRN=8'hB8;
            BLU=8'h88;
        end
        1942:
        begin
            RED=8'hBE;
            GRN=8'hCC;
            BLU=8'hBA;
        end
        1943:
        begin
            RED=8'hB9;
            GRN=8'hD8;
            BLU=8'hD2;
        end
        1944:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1945:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1946:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1947:
        begin
            RED=8'hB7;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        1948:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        1949:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        1950:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        1951:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        1952:
        begin
            RED=8'hB5;
            GRN=8'hD7;
            BLU=8'hD0;
        end
        1953:
        begin
            RED=8'h91;
            GRN=8'hB9;
            BLU=8'hB1;
        end
        1954:
        begin
            RED=8'h8B;
            GRN=8'hBC;
            BLU=8'hB3;
        end
        1955:
        begin
            RED=8'h8E;
            GRN=8'hC3;
            BLU=8'hBB;
        end
        1956:
        begin
            RED=8'h8E;
            GRN=8'hC2;
            BLU=8'hBD;
        end
        1957:
        begin
            RED=8'h91;
            GRN=8'hC0;
            BLU=8'hBB;
        end
        1958:
        begin
            RED=8'h9E;
            GRN=8'hAD;
            BLU=8'h94;
        end
        1959:
        begin
            RED=8'hE0;
            GRN=8'hBF;
            BLU=8'h86;
        end
        1960:
        begin
            RED=8'hF1;
            GRN=8'hC1;
            BLU=8'h7F;
        end
        1961:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1962:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        1963:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h81;
        end
        1964:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h84;
        end
        1965:
        begin
            RED=8'hEB;
            GRN=8'hC0;
            BLU=8'h84;
        end
        1966:
        begin
            RED=8'hE8;
            GRN=8'hC0;
            BLU=8'h88;
        end
        1967:
        begin
            RED=8'hE5;
            GRN=8'hBD;
            BLU=8'h85;
        end
        1968:
        begin
            RED=8'hDE;
            GRN=8'hB7;
            BLU=8'h7E;
        end
        1969:
        begin
            RED=8'hD5;
            GRN=8'hAE;
            BLU=8'h75;
        end
        1970:
        begin
            RED=8'hAF;
            GRN=8'h96;
            BLU=8'h66;
        end
        1971:
        begin
            RED=8'h74;
            GRN=8'h6B;
            BLU=8'h47;
        end
        1972:
        begin
            RED=8'h75;
            GRN=8'h7A;
            BLU=8'h5F;
        end
        1973:
        begin
            RED=8'h7D;
            GRN=8'h85;
            BLU=8'h67;
        end
        1974:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h61;
        end
        1975:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        1976:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        1977:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h68;
        end
        1978:
        begin
            RED=8'h55;
            GRN=8'h57;
            BLU=8'h49;
        end
        1979:
        begin
            RED=8'h2E;
            GRN=8'h2F;
            BLU=8'h27;
        end
        1980:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1981:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1982:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1983:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        1984:
        begin
            RED=8'h7A;
            GRN=8'h85;
            BLU=8'h65;
        end
        1985:
        begin
            RED=8'h7E;
            GRN=8'h84;
            BLU=8'h62;
        end
        1986:
        begin
            RED=8'h81;
            GRN=8'h83;
            BLU=8'h60;
        end
        1987:
        begin
            RED=8'h81;
            GRN=8'h83;
            BLU=8'h64;
        end
        1988:
        begin
            RED=8'h7A;
            GRN=8'h80;
            BLU=8'h67;
        end
        1989:
        begin
            RED=8'h6D;
            GRN=8'h7C;
            BLU=8'h6E;
        end
        1990:
        begin
            RED=8'hA9;
            GRN=8'hCA;
            BLU=8'hBB;
        end
        1991:
        begin
            RED=8'hB4;
            GRN=8'hDB;
            BLU=8'hD0;
        end
        1992:
        begin
            RED=8'hB9;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        1993:
        begin
            RED=8'hB8;
            GRN=8'hD9;
            BLU=8'hD1;
        end
        1994:
        begin
            RED=8'hB4;
            GRN=8'hDA;
            BLU=8'hD3;
        end
        1995:
        begin
            RED=8'hB6;
            GRN=8'hD7;
            BLU=8'hD4;
        end
        1996:
        begin
            RED=8'hC4;
            GRN=8'hD1;
            BLU=8'hC5;
        end
        1997:
        begin
            RED=8'hB4;
            GRN=8'hA9;
            BLU=8'h8C;
        end
        1998:
        begin
            RED=8'hEB;
            GRN=8'hBF;
            BLU=8'h84;
        end
        1999:
        begin
            RED=8'hED;
            GRN=8'hBD;
            BLU=8'h82;
        end
        2000:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h81;
        end
        2001:
        begin
            RED=8'hEB;
            GRN=8'hC1;
            BLU=8'h7F;
        end
        2002:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        2003:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h84;
        end
        2004:
        begin
            RED=8'hEB;
            GRN=8'hC1;
            BLU=8'h7A;
        end
        2005:
        begin
            RED=8'hEC;
            GRN=8'hC1;
            BLU=8'h7D;
        end
        2006:
        begin
            RED=8'hBB;
            GRN=8'hB4;
            BLU=8'h94;
        end
        2007:
        begin
            RED=8'hB8;
            GRN=8'hD4;
            BLU=8'hCD;
        end
        2008:
        begin
            RED=8'hB5;
            GRN=8'hD5;
            BLU=8'hD0;
        end
        2009:
        begin
            RED=8'hB8;
            GRN=8'hD9;
            BLU=8'hD4;
        end
        2010:
        begin
            RED=8'hB8;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        2011:
        begin
            RED=8'hB7;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        2012:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        2013:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        2014:
        begin
            RED=8'hB6;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        2015:
        begin
            RED=8'hB7;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        2016:
        begin
            RED=8'hA8;
            GRN=8'hC8;
            BLU=8'hC2;
        end
        2017:
        begin
            RED=8'h7F;
            GRN=8'hAB;
            BLU=8'hA2;
        end
        2018:
        begin
            RED=8'h8C;
            GRN=8'hC3;
            BLU=8'hB8;
        end
        2019:
        begin
            RED=8'h8D;
            GRN=8'hC3;
            BLU=8'hBB;
        end
        2020:
        begin
            RED=8'h91;
            GRN=8'hC2;
            BLU=8'hBC;
        end
        2021:
        begin
            RED=8'h99;
            GRN=8'hBD;
            BLU=8'hB5;
        end
        2022:
        begin
            RED=8'h9C;
            GRN=8'h9B;
            BLU=8'h7B;
        end
        2023:
        begin
            RED=8'hE8;
            GRN=8'hC0;
            BLU=8'h82;
        end
        2024:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h80;
        end
        2025:
        begin
            RED=8'hEC;
            GRN=8'hC1;
            BLU=8'h7D;
        end
        2026:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7C;
        end
        2027:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        2028:
        begin
            RED=8'hEC;
            GRN=8'hBE;
            BLU=8'h80;
        end
        2029:
        begin
            RED=8'hE4;
            GRN=8'hB7;
            BLU=8'h7C;
        end
        2030:
        begin
            RED=8'hC6;
            GRN=8'h9F;
            BLU=8'h6A;
        end
        2031:
        begin
            RED=8'hC3;
            GRN=8'h9C;
            BLU=8'h67;
        end
        2032:
        begin
            RED=8'hCE;
            GRN=8'hA7;
            BLU=8'h73;
        end
        2033:
        begin
            RED=8'hC6;
            GRN=8'h9F;
            BLU=8'h6A;
        end
        2034:
        begin
            RED=8'h8C;
            GRN=8'h7A;
            BLU=8'h52;
        end
        2035:
        begin
            RED=8'h7D;
            GRN=8'h7F;
            BLU=8'h62;
        end
        2036:
        begin
            RED=8'h69;
            GRN=8'h75;
            BLU=8'h5E;
        end
        2037:
        begin
            RED=8'h65;
            GRN=8'h6E;
            BLU=8'h51;
        end
        2038:
        begin
            RED=8'h80;
            GRN=8'h82;
            BLU=8'h61;
        end
        2039:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        2040:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2041:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h68;
        end
        2042:
        begin
            RED=8'h55;
            GRN=8'h57;
            BLU=8'h49;
        end
        2043:
        begin
            RED=8'h2E;
            GRN=8'h2F;
            BLU=8'h27;
        end
        2044:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2045:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2046:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2047:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2048:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2049:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2050:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2051:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2052:
        begin
            RED=8'h7E;
            GRN=8'h84;
            BLU=8'h66;
        end
        2053:
        begin
            RED=8'h78;
            GRN=8'h84;
            BLU=8'h6B;
        end
        2054:
        begin
            RED=8'h72;
            GRN=8'h86;
            BLU=8'h73;
        end
        2055:
        begin
            RED=8'h8B;
            GRN=8'hA4;
            BLU=8'h97;
        end
        2056:
        begin
            RED=8'hB6;
            GRN=8'hCF;
            BLU=8'hC5;
        end
        2057:
        begin
            RED=8'hBC;
            GRN=8'hD7;
            BLU=8'hD2;
        end
        2058:
        begin
            RED=8'hB6;
            GRN=8'hD8;
            BLU=8'hCC;
        end
        2059:
        begin
            RED=8'hB9;
            GRN=8'hD1;
            BLU=8'hC6;
        end
        2060:
        begin
            RED=8'hAB;
            GRN=8'hA2;
            BLU=8'h8B;
        end
        2061:
        begin
            RED=8'hE3;
            GRN=8'hBD;
            BLU=8'h87;
        end
        2062:
        begin
            RED=8'hEF;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2063:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h7F;
        end
        2064:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2065:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2066:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2067:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2068:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2069:
        begin
            RED=8'hEA;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2070:
        begin
            RED=8'hE2;
            GRN=8'hC0;
            BLU=8'h8A;
        end
        2071:
        begin
            RED=8'hB1;
            GRN=8'hAB;
            BLU=8'h92;
        end
        2072:
        begin
            RED=8'hB4;
            GRN=8'hC8;
            BLU=8'hB8;
        end
        2073:
        begin
            RED=8'hB5;
            GRN=8'hDB;
            BLU=8'hD1;
        end
        2074:
        begin
            RED=8'hB7;
            GRN=8'hDA;
            BLU=8'hD5;
        end
        2075:
        begin
            RED=8'hB9;
            GRN=8'hD8;
            BLU=8'hD3;
        end
        2076:
        begin
            RED=8'hB8;
            GRN=8'hD9;
            BLU=8'hD3;
        end
        2077:
        begin
            RED=8'hB7;
            GRN=8'hD9;
            BLU=8'hD2;
        end
        2078:
        begin
            RED=8'hB5;
            GRN=8'hD8;
            BLU=8'hCF;
        end
        2079:
        begin
            RED=8'h9A;
            GRN=8'hBE;
            BLU=8'hB4;
        end
        2080:
        begin
            RED=8'h83;
            GRN=8'hAA;
            BLU=8'hA2;
        end
        2081:
        begin
            RED=8'h91;
            GRN=8'hC1;
            BLU=8'hBB;
        end
        2082:
        begin
            RED=8'h8E;
            GRN=8'hC3;
            BLU=8'hBD;
        end
        2083:
        begin
            RED=8'h91;
            GRN=8'hC5;
            BLU=8'hBC;
        end
        2084:
        begin
            RED=8'h97;
            GRN=8'hC1;
            BLU=8'hB2;
        end
        2085:
        begin
            RED=8'h9A;
            GRN=8'hA5;
            BLU=8'h88;
        end
        2086:
        begin
            RED=8'hD9;
            GRN=8'hBD;
            BLU=8'h8E;
        end
        2087:
        begin
            RED=8'hF0;
            GRN=8'hBF;
            BLU=8'h7F;
        end
        2088:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h7C;
        end
        2089:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        2090:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        2091:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        2092:
        begin
            RED=8'hE3;
            GRN=8'hB6;
            BLU=8'h75;
        end
        2093:
        begin
            RED=8'hD5;
            GRN=8'hA8;
            BLU=8'h6B;
        end
        2094:
        begin
            RED=8'hE7;
            GRN=8'hBD;
            BLU=8'h83;
        end
        2095:
        begin
            RED=8'hE9;
            GRN=8'hC0;
            BLU=8'h83;
        end
        2096:
        begin
            RED=8'hE7;
            GRN=8'hBF;
            BLU=8'h8A;
        end
        2097:
        begin
            RED=8'hE8;
            GRN=8'hC3;
            BLU=8'h84;
        end
        2098:
        begin
            RED=8'hDE;
            GRN=8'hBD;
            BLU=8'h80;
        end
        2099:
        begin
            RED=8'h84;
            GRN=8'h7E;
            BLU=8'h5D;
        end
        2100:
        begin
            RED=8'h76;
            GRN=8'h85;
            BLU=8'h70;
        end
        2101:
        begin
            RED=8'h6D;
            GRN=8'h75;
            BLU=8'h57;
        end
        2102:
        begin
            RED=8'h7D;
            GRN=8'h80;
            BLU=8'h5F;
        end
        2103:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        2104:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2105:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h69;
        end
        2106:
        begin
            RED=8'h56;
            GRN=8'h58;
            BLU=8'h4A;
        end
        2107:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h28;
        end
        2108:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2109:
        begin
            RED=8'h31;
            GRN=8'h32;
            BLU=8'h2A;
        end
        2110:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2111:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2112:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2113:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2114:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2115:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2116:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h62;
        end
        2117:
        begin
            RED=8'h81;
            GRN=8'h83;
            BLU=8'h5F;
        end
        2118:
        begin
            RED=8'h80;
            GRN=8'h81;
            BLU=8'h60;
        end
        2119:
        begin
            RED=8'h83;
            GRN=8'h7D;
            BLU=8'h5A;
        end
        2120:
        begin
            RED=8'hC7;
            GRN=8'hB8;
            BLU=8'h8D;
        end
        2121:
        begin
            RED=8'hBC;
            GRN=8'hA9;
            BLU=8'h81;
        end
        2122:
        begin
            RED=8'hB2;
            GRN=8'hA6;
            BLU=8'h7B;
        end
        2123:
        begin
            RED=8'hBB;
            GRN=8'hAF;
            BLU=8'h89;
        end
        2124:
        begin
            RED=8'hB7;
            GRN=8'h98;
            BLU=8'h6E;
        end
        2125:
        begin
            RED=8'hEF;
            GRN=8'hC1;
            BLU=8'h7D;
        end
        2126:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2127:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2128:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2129:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2130:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2131:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2132:
        begin
            RED=8'hEB;
            GRN=8'hC0;
            BLU=8'h81;
        end
        2133:
        begin
            RED=8'hE9;
            GRN=8'hC0;
            BLU=8'h82;
        end
        2134:
        begin
            RED=8'hE9;
            GRN=8'hC1;
            BLU=8'h84;
        end
        2135:
        begin
            RED=8'hE8;
            GRN=8'hC2;
            BLU=8'h82;
        end
        2136:
        begin
            RED=8'hD0;
            GRN=8'hB7;
            BLU=8'h86;
        end
        2137:
        begin
            RED=8'hAA;
            GRN=8'hA6;
            BLU=8'h8A;
        end
        2138:
        begin
            RED=8'hB3;
            GRN=8'hC2;
            BLU=8'hB2;
        end
        2139:
        begin
            RED=8'hB2;
            GRN=8'hCD;
            BLU=8'hBF;
        end
        2140:
        begin
            RED=8'hAB;
            GRN=8'hCC;
            BLU=8'hBD;
        end
        2141:
        begin
            RED=8'h9E;
            GRN=8'hC4;
            BLU=8'hB7;
        end
        2142:
        begin
            RED=8'h87;
            GRN=8'hB2;
            BLU=8'hA6;
        end
        2143:
        begin
            RED=8'h8B;
            GRN=8'hBB;
            BLU=8'hB0;
        end
        2144:
        begin
            RED=8'h8B;
            GRN=8'hC3;
            BLU=8'hB9;
        end
        2145:
        begin
            RED=8'h8A;
            GRN=8'hC5;
            BLU=8'hBC;
        end
        2146:
        begin
            RED=8'h8D;
            GRN=8'hC3;
            BLU=8'hB9;
        end
        2147:
        begin
            RED=8'h93;
            GRN=8'hBF;
            BLU=8'hAE;
        end
        2148:
        begin
            RED=8'h91;
            GRN=8'hA9;
            BLU=8'h8D;
        end
        2149:
        begin
            RED=8'hC3;
            GRN=8'hB5;
            BLU=8'h86;
        end
        2150:
        begin
            RED=8'hEC;
            GRN=8'hC2;
            BLU=8'h88;
        end
        2151:
        begin
            RED=8'hF1;
            GRN=8'hBE;
            BLU=8'h7D;
        end
        2152:
        begin
            RED=8'hE9;
            GRN=8'hC2;
            BLU=8'h7E;
        end
        2153:
        begin
            RED=8'hEB;
            GRN=8'hC1;
            BLU=8'h7F;
        end
        2154:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2155:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2156:
        begin
            RED=8'hEE;
            GRN=8'hC1;
            BLU=8'h80;
        end
        2157:
        begin
            RED=8'hEC;
            GRN=8'hBE;
            BLU=8'h81;
        end
        2158:
        begin
            RED=8'hDF;
            GRN=8'hB3;
            BLU=8'h7E;
        end
        2159:
        begin
            RED=8'hC2;
            GRN=8'h98;
            BLU=8'h65;
        end
        2160:
        begin
            RED=8'hA1;
            GRN=8'h75;
            BLU=8'h56;
        end
        2161:
        begin
            RED=8'hC2;
            GRN=8'h99;
            BLU=8'h6E;
        end
        2162:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h83;
        end
        2163:
        begin
            RED=8'hAA;
            GRN=8'h9C;
            BLU=8'h74;
        end
        2164:
        begin
            RED=8'h79;
            GRN=8'h83;
            BLU=8'h6A;
        end
        2165:
        begin
            RED=8'h7E;
            GRN=8'h84;
            BLU=8'h66;
        end
        2166:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h64;
        end
        2167:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        2168:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2169:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h69;
        end
        2170:
        begin
            RED=8'h56;
            GRN=8'h58;
            BLU=8'h4A;
        end
        2171:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h28;
        end
        2172:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2173:
        begin
            RED=8'h31;
            GRN=8'h32;
            BLU=8'h2A;
        end
        2174:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2175:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2176:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2177:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2178:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2179:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2180:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h62;
        end
        2181:
        begin
            RED=8'h7D;
            GRN=8'h82;
            BLU=8'h61;
        end
        2182:
        begin
            RED=8'h81;
            GRN=8'h83;
            BLU=8'h63;
        end
        2183:
        begin
            RED=8'h89;
            GRN=8'h7B;
            BLU=8'h52;
        end
        2184:
        begin
            RED=8'hE2;
            GRN=8'hBE;
            BLU=8'h83;
        end
        2185:
        begin
            RED=8'hED;
            GRN=8'hBE;
            BLU=8'h83;
        end
        2186:
        begin
            RED=8'hDF;
            GRN=8'hB9;
            BLU=8'h7B;
        end
        2187:
        begin
            RED=8'hC9;
            GRN=8'hAA;
            BLU=8'h75;
        end
        2188:
        begin
            RED=8'hD0;
            GRN=8'hAB;
            BLU=8'h7A;
        end
        2189:
        begin
            RED=8'hE9;
            GRN=8'hBF;
            BLU=8'h7C;
        end
        2190:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2191:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2192:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2193:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2194:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2195:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2196:
        begin
            RED=8'hE7;
            GRN=8'hBC;
            BLU=8'h7D;
        end
        2197:
        begin
            RED=8'hCD;
            GRN=8'hA5;
            BLU=8'h67;
        end
        2198:
        begin
            RED=8'hD3;
            GRN=8'hAB;
            BLU=8'h6D;
        end
        2199:
        begin
            RED=8'hE6;
            GRN=8'hC1;
            BLU=8'h78;
        end
        2200:
        begin
            RED=8'hF0;
            GRN=8'hBE;
            BLU=8'h7E;
        end
        2201:
        begin
            RED=8'hEF;
            GRN=8'hBC;
            BLU=8'h87;
        end
        2202:
        begin
            RED=8'hDC;
            GRN=8'hBA;
            BLU=8'h8A;
        end
        2203:
        begin
            RED=8'hB9;
            GRN=8'hA6;
            BLU=8'h7A;
        end
        2204:
        begin
            RED=8'hA8;
            GRN=8'h9C;
            BLU=8'h77;
        end
        2205:
        begin
            RED=8'hA0;
            GRN=8'h9A;
            BLU=8'h78;
        end
        2206:
        begin
            RED=8'h9F;
            GRN=8'hA2;
            BLU=8'h84;
        end
        2207:
        begin
            RED=8'hA1;
            GRN=8'hAB;
            BLU=8'h90;
        end
        2208:
        begin
            RED=8'hA0;
            GRN=8'hB0;
            BLU=8'h92;
        end
        2209:
        begin
            RED=8'hA0;
            GRN=8'hAE;
            BLU=8'h91;
        end
        2210:
        begin
            RED=8'hA3;
            GRN=8'hA8;
            BLU=8'h87;
        end
        2211:
        begin
            RED=8'hAE;
            GRN=8'hA3;
            BLU=8'h7B;
        end
        2212:
        begin
            RED=8'hD7;
            GRN=8'hBE;
            BLU=8'h8C;
        end
        2213:
        begin
            RED=8'hE9;
            GRN=8'hC3;
            BLU=8'h83;
        end
        2214:
        begin
            RED=8'hF1;
            GRN=8'hC1;
            BLU=8'h7F;
        end
        2215:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h7C;
        end
        2216:
        begin
            RED=8'hE9;
            GRN=8'hC2;
            BLU=8'h80;
        end
        2217:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2218:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2219:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2220:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        2221:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h7F;
        end
        2222:
        begin
            RED=8'hE0;
            GRN=8'hB6;
            BLU=8'h75;
        end
        2223:
        begin
            RED=8'hE9;
            GRN=8'hC0;
            BLU=8'h84;
        end
        2224:
        begin
            RED=8'hDD;
            GRN=8'hB1;
            BLU=8'h89;
        end
        2225:
        begin
            RED=8'hCB;
            GRN=8'hA3;
            BLU=8'h75;
        end
        2226:
        begin
            RED=8'hE7;
            GRN=8'hC0;
            BLU=8'h84;
        end
        2227:
        begin
            RED=8'h98;
            GRN=8'h8A;
            BLU=8'h61;
        end
        2228:
        begin
            RED=8'h7D;
            GRN=8'h82;
            BLU=8'h65;
        end
        2229:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h63;
        end
        2230:
        begin
            RED=8'h7A;
            GRN=8'h83;
            BLU=8'h65;
        end
        2231:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        2232:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2233:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h69;
        end
        2234:
        begin
            RED=8'h56;
            GRN=8'h58;
            BLU=8'h4A;
        end
        2235:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h28;
        end
        2236:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2237:
        begin
            RED=8'h31;
            GRN=8'h32;
            BLU=8'h2A;
        end
        2238:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2239:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2240:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2241:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2242:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2243:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2244:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h62;
        end
        2245:
        begin
            RED=8'h7D;
            GRN=8'h83;
            BLU=8'h65;
        end
        2246:
        begin
            RED=8'h78;
            GRN=8'h84;
            BLU=8'h6B;
        end
        2247:
        begin
            RED=8'h80;
            GRN=8'h7F;
            BLU=8'h5F;
        end
        2248:
        begin
            RED=8'hA4;
            GRN=8'h8A;
            BLU=8'h58;
        end
        2249:
        begin
            RED=8'hE3;
            GRN=8'hBA;
            BLU=8'h87;
        end
        2250:
        begin
            RED=8'hC6;
            GRN=8'hA1;
            BLU=8'h65;
        end
        2251:
        begin
            RED=8'hDA;
            GRN=8'hB8;
            BLU=8'h80;
        end
        2252:
        begin
            RED=8'hDD;
            GRN=8'hB7;
            BLU=8'h82;
        end
        2253:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h7D;
        end
        2254:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2255:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2256:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2257:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2258:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2259:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2260:
        begin
            RED=8'hEB;
            GRN=8'hC0;
            BLU=8'h81;
        end
        2261:
        begin
            RED=8'hEB;
            GRN=8'hC3;
            BLU=8'h85;
        end
        2262:
        begin
            RED=8'hD9;
            GRN=8'hB1;
            BLU=8'h75;
        end
        2263:
        begin
            RED=8'hDD;
            GRN=8'hB8;
            BLU=8'h83;
        end
        2264:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h84;
        end
        2265:
        begin
            RED=8'hF1;
            GRN=8'hBD;
            BLU=8'h7C;
        end
        2266:
        begin
            RED=8'hF2;
            GRN=8'hBE;
            BLU=8'h7D;
        end
        2267:
        begin
            RED=8'hEF;
            GRN=8'hBE;
            BLU=8'h82;
        end
        2268:
        begin
            RED=8'hE8;
            GRN=8'hB9;
            BLU=8'h83;
        end
        2269:
        begin
            RED=8'hC5;
            GRN=8'h9A;
            BLU=8'h65;
        end
        2270:
        begin
            RED=8'hE4;
            GRN=8'hBE;
            BLU=8'h88;
        end
        2271:
        begin
            RED=8'hE4;
            GRN=8'hC1;
            BLU=8'h8C;
        end
        2272:
        begin
            RED=8'hE5;
            GRN=8'hBF;
            BLU=8'h88;
        end
        2273:
        begin
            RED=8'hE5;
            GRN=8'hC0;
            BLU=8'h8A;
        end
        2274:
        begin
            RED=8'hE6;
            GRN=8'hBF;
            BLU=8'h87;
        end
        2275:
        begin
            RED=8'hEF;
            GRN=8'hC1;
            BLU=8'h83;
        end
        2276:
        begin
            RED=8'hF1;
            GRN=8'hBF;
            BLU=8'h7C;
        end
        2277:
        begin
            RED=8'hEF;
            GRN=8'hC1;
            BLU=8'h7D;
        end
        2278:
        begin
            RED=8'hEE;
            GRN=8'hC2;
            BLU=8'h7E;
        end
        2279:
        begin
            RED=8'hEB;
            GRN=8'hC1;
            BLU=8'h7E;
        end
        2280:
        begin
            RED=8'hEB;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2281:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2282:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2283:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2284:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2285:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2286:
        begin
            RED=8'hEC;
            GRN=8'hC3;
            BLU=8'h7F;
        end
        2287:
        begin
            RED=8'hE9;
            GRN=8'hC1;
            BLU=8'h7E;
        end
        2288:
        begin
            RED=8'hCD;
            GRN=8'hA4;
            BLU=8'h6F;
        end
        2289:
        begin
            RED=8'hE6;
            GRN=8'hC0;
            BLU=8'h83;
        end
        2290:
        begin
            RED=8'hD6;
            GRN=8'hBB;
            BLU=8'h83;
        end
        2291:
        begin
            RED=8'h7A;
            GRN=8'h77;
            BLU=8'h57;
        end
        2292:
        begin
            RED=8'h7D;
            GRN=8'h85;
            BLU=8'h6B;
        end
        2293:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h63;
        end
        2294:
        begin
            RED=8'h7C;
            GRN=8'h84;
            BLU=8'h66;
        end
        2295:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        2296:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2297:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h69;
        end
        2298:
        begin
            RED=8'h55;
            GRN=8'h57;
            BLU=8'h4A;
        end
        2299:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h28;
        end
        2300:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2301:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2302:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2303:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2304:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2305:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2306:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2307:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2308:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h61;
        end
        2309:
        begin
            RED=8'h81;
            GRN=8'h82;
            BLU=8'h5E;
        end
        2310:
        begin
            RED=8'h7C;
            GRN=8'h83;
            BLU=8'h69;
        end
        2311:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h65;
        end
        2312:
        begin
            RED=8'hA3;
            GRN=8'h8F;
            BLU=8'h62;
        end
        2313:
        begin
            RED=8'hD3;
            GRN=8'hAD;
            BLU=8'h7D;
        end
        2314:
        begin
            RED=8'hD5;
            GRN=8'hB0;
            BLU=8'h7A;
        end
        2315:
        begin
            RED=8'hCE;
            GRN=8'hAA;
            BLU=8'h72;
        end
        2316:
        begin
            RED=8'hE4;
            GRN=8'hBA;
            BLU=8'h7E;
        end
        2317:
        begin
            RED=8'hEF;
            GRN=8'hC1;
            BLU=8'h76;
        end
        2318:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2319:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2320:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2321:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        2322:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2323:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2324:
        begin
            RED=8'hEA;
            GRN=8'hC0;
            BLU=8'h82;
        end
        2325:
        begin
            RED=8'hE8;
            GRN=8'hC0;
            BLU=8'h84;
        end
        2326:
        begin
            RED=8'hDB;
            GRN=8'hB2;
            BLU=8'h79;
        end
        2327:
        begin
            RED=8'hE4;
            GRN=8'hB3;
            BLU=8'h7E;
        end
        2328:
        begin
            RED=8'hEC;
            GRN=8'hC1;
            BLU=8'h83;
        end
        2329:
        begin
            RED=8'hEA;
            GRN=8'hC3;
            BLU=8'h82;
        end
        2330:
        begin
            RED=8'hD9;
            GRN=8'hB0;
            BLU=8'h7A;
        end
        2331:
        begin
            RED=8'hE5;
            GRN=8'hBB;
            BLU=8'h86;
        end
        2332:
        begin
            RED=8'hEA;
            GRN=8'hC2;
            BLU=8'h83;
        end
        2333:
        begin
            RED=8'hE0;
            GRN=8'hB8;
            BLU=8'h77;
        end
        2334:
        begin
            RED=8'hC6;
            GRN=8'h9E;
            BLU=8'h5F;
        end
        2335:
        begin
            RED=8'hDB;
            GRN=8'hB3;
            BLU=8'h77;
        end
        2336:
        begin
            RED=8'hEE;
            GRN=8'hBE;
            BLU=8'h7E;
        end
        2337:
        begin
            RED=8'hEF;
            GRN=8'hC1;
            BLU=8'h82;
        end
        2338:
        begin
            RED=8'hEC;
            GRN=8'hC4;
            BLU=8'h84;
        end
        2339:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h7F;
        end
        2340:
        begin
            RED=8'hEB;
            GRN=8'hBF;
            BLU=8'h7B;
        end
        2341:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        2342:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h80;
        end
        2343:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h7F;
        end
        2344:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2345:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2346:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2347:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2348:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        2349:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2350:
        begin
            RED=8'hE8;
            GRN=8'hBF;
            BLU=8'h87;
        end
        2351:
        begin
            RED=8'hDA;
            GRN=8'hAE;
            BLU=8'h74;
        end
        2352:
        begin
            RED=8'hD3;
            GRN=8'hAA;
            BLU=8'h6E;
        end
        2353:
        begin
            RED=8'hE2;
            GRN=8'hC3;
            BLU=8'h86;
        end
        2354:
        begin
            RED=8'h8F;
            GRN=8'h84;
            BLU=8'h58;
        end
        2355:
        begin
            RED=8'h7B;
            GRN=8'h81;
            BLU=8'h66;
        end
        2356:
        begin
            RED=8'h7B;
            GRN=8'h84;
            BLU=8'h69;
        end
        2357:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h62;
        end
        2358:
        begin
            RED=8'h7C;
            GRN=8'h84;
            BLU=8'h65;
        end
        2359:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        2360:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2361:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h69;
        end
        2362:
        begin
            RED=8'h54;
            GRN=8'h59;
            BLU=8'h4A;
        end
        2363:
        begin
            RED=8'h2F;
            GRN=8'h31;
            BLU=8'h29;
        end
        2364:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2365:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2366:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2367:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2368:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2369:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2370:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2371:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2372:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h63;
        end
        2373:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h63;
        end
        2374:
        begin
            RED=8'h7F;
            GRN=8'h81;
            BLU=8'h69;
        end
        2375:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2376:
        begin
            RED=8'h9E;
            GRN=8'h8D;
            BLU=8'h62;
        end
        2377:
        begin
            RED=8'hE6;
            GRN=8'hBE;
            BLU=8'h88;
        end
        2378:
        begin
            RED=8'hC1;
            GRN=8'h9A;
            BLU=8'h65;
        end
        2379:
        begin
            RED=8'hD1;
            GRN=8'hAF;
            BLU=8'h7D;
        end
        2380:
        begin
            RED=8'hE7;
            GRN=8'hC1;
            BLU=8'h85;
        end
        2381:
        begin
            RED=8'hEE;
            GRN=8'hC3;
            BLU=8'h7C;
        end
        2382:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2383:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2384:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h82;
        end
        2385:
        begin
            RED=8'hEE;
            GRN=8'hC1;
            BLU=8'h84;
        end
        2386:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h83;
        end
        2387:
        begin
            RED=8'hE8;
            GRN=8'hBE;
            BLU=8'h82;
        end
        2388:
        begin
            RED=8'hE9;
            GRN=8'hC0;
            BLU=8'h85;
        end
        2389:
        begin
            RED=8'hE1;
            GRN=8'hBA;
            BLU=8'h80;
        end
        2390:
        begin
            RED=8'hC7;
            GRN=8'hA2;
            BLU=8'h67;
        end
        2391:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h80;
        end
        2392:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        2393:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        2394:
        begin
            RED=8'hEA;
            GRN=8'hBB;
            BLU=8'h87;
        end
        2395:
        begin
            RED=8'hD5;
            GRN=8'hA8;
            BLU=8'h73;
        end
        2396:
        begin
            RED=8'hE9;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        2397:
        begin
            RED=8'hEB;
            GRN=8'hC3;
            BLU=8'h7C;
        end
        2398:
        begin
            RED=8'hE9;
            GRN=8'hC1;
            BLU=8'h7F;
        end
        2399:
        begin
            RED=8'hDE;
            GRN=8'hB3;
            BLU=8'h7B;
        end
        2400:
        begin
            RED=8'hD3;
            GRN=8'hA5;
            BLU=8'h69;
        end
        2401:
        begin
            RED=8'hCC;
            GRN=8'h9E;
            BLU=8'h60;
        end
        2402:
        begin
            RED=8'hD8;
            GRN=8'hAA;
            BLU=8'h6C;
        end
        2403:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h82;
        end
        2404:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h81;
        end
        2405:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2406:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2407:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2408:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2409:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        2410:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2411:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2412:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        2413:
        begin
            RED=8'hEB;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2414:
        begin
            RED=8'hCA;
            GRN=8'hA2;
            BLU=8'h6E;
        end
        2415:
        begin
            RED=8'hDD;
            GRN=8'hAC;
            BLU=8'h71;
        end
        2416:
        begin
            RED=8'hE8;
            GRN=8'hC2;
            BLU=8'h80;
        end
        2417:
        begin
            RED=8'h9B;
            GRN=8'h8E;
            BLU=8'h61;
        end
        2418:
        begin
            RED=8'h7B;
            GRN=8'h7D;
            BLU=8'h5D;
        end
        2419:
        begin
            RED=8'h7D;
            GRN=8'h82;
            BLU=8'h62;
        end
        2420:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2421:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2422:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2423:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        2424:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h63;
        end
        2425:
        begin
            RED=8'h7C;
            GRN=8'h85;
            BLU=8'h6A;
        end
        2426:
        begin
            RED=8'h53;
            GRN=8'h5B;
            BLU=8'h4B;
        end
        2427:
        begin
            RED=8'h2F;
            GRN=8'h33;
            BLU=8'h29;
        end
        2428:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2429:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2430:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2431:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2432:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2433:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2434:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2435:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2436:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h63;
        end
        2437:
        begin
            RED=8'h7C;
            GRN=8'h84;
            BLU=8'h63;
        end
        2438:
        begin
            RED=8'h80;
            GRN=8'h81;
            BLU=8'h67;
        end
        2439:
        begin
            RED=8'h7A;
            GRN=8'h83;
            BLU=8'h61;
        end
        2440:
        begin
            RED=8'h83;
            GRN=8'h7C;
            BLU=8'h54;
        end
        2441:
        begin
            RED=8'hDE;
            GRN=8'hBD;
            BLU=8'h85;
        end
        2442:
        begin
            RED=8'hDC;
            GRN=8'hB6;
            BLU=8'h7C;
        end
        2443:
        begin
            RED=8'hDC;
            GRN=8'hB3;
            BLU=8'h7E;
        end
        2444:
        begin
            RED=8'hEB;
            GRN=8'hBF;
            BLU=8'h85;
        end
        2445:
        begin
            RED=8'hEC;
            GRN=8'hBD;
            BLU=8'h7C;
        end
        2446:
        begin
            RED=8'hEB;
            GRN=8'hC1;
            BLU=8'h7D;
        end
        2447:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2448:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h84;
        end
        2449:
        begin
            RED=8'hDF;
            GRN=8'hB2;
            BLU=8'h7B;
        end
        2450:
        begin
            RED=8'hCB;
            GRN=8'h9D;
            BLU=8'h67;
        end
        2451:
        begin
            RED=8'hC7;
            GRN=8'h9A;
            BLU=8'h62;
        end
        2452:
        begin
            RED=8'hCB;
            GRN=8'hA1;
            BLU=8'h66;
        end
        2453:
        begin
            RED=8'hD4;
            GRN=8'hAD;
            BLU=8'h6D;
        end
        2454:
        begin
            RED=8'hE8;
            GRN=8'hC1;
            BLU=8'h7F;
        end
        2455:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2456:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2457:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h80;
        end
        2458:
        begin
            RED=8'hED;
            GRN=8'hBE;
            BLU=8'h86;
        end
        2459:
        begin
            RED=8'hD2;
            GRN=8'hA5;
            BLU=8'h71;
        end
        2460:
        begin
            RED=8'hE8;
            GRN=8'hBD;
            BLU=8'h86;
        end
        2461:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h83;
        end
        2462:
        begin
            RED=8'hE8;
            GRN=8'hBF;
            BLU=8'h7C;
        end
        2463:
        begin
            RED=8'hE9;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        2464:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h80;
        end
        2465:
        begin
            RED=8'hEF;
            GRN=8'hC1;
            BLU=8'h81;
        end
        2466:
        begin
            RED=8'hEC;
            GRN=8'hBE;
            BLU=8'h7E;
        end
        2467:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2468:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2469:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2470:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2471:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2472:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2473:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2474:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2475:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h80;
        end
        2476:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        2477:
        begin
            RED=8'hE8;
            GRN=8'hBA;
            BLU=8'h82;
        end
        2478:
        begin
            RED=8'hD1;
            GRN=8'hA4;
            BLU=8'h70;
        end
        2479:
        begin
            RED=8'hE9;
            GRN=8'hC1;
            BLU=8'h82;
        end
        2480:
        begin
            RED=8'hBF;
            GRN=8'hA5;
            BLU=8'h82;
        end
        2481:
        begin
            RED=8'h7B;
            GRN=8'h79;
            BLU=8'h5B;
        end
        2482:
        begin
            RED=8'h80;
            GRN=8'h86;
            BLU=8'h64;
        end
        2483:
        begin
            RED=8'h7F;
            GRN=8'h84;
            BLU=8'h64;
        end
        2484:
        begin
            RED=8'h7D;
            GRN=8'h82;
            BLU=8'h62;
        end
        2485:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2486:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2487:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        2488:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h63;
        end
        2489:
        begin
            RED=8'h7C;
            GRN=8'h85;
            BLU=8'h6A;
        end
        2490:
        begin
            RED=8'h53;
            GRN=8'h5B;
            BLU=8'h4B;
        end
        2491:
        begin
            RED=8'h2F;
            GRN=8'h33;
            BLU=8'h29;
        end
        2492:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2493:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2494:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2495:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2496:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2497:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2498:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2499:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2500:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h63;
        end
        2501:
        begin
            RED=8'h7C;
            GRN=8'h84;
            BLU=8'h65;
        end
        2502:
        begin
            RED=8'h81;
            GRN=8'h82;
            BLU=8'h64;
        end
        2503:
        begin
            RED=8'h7A;
            GRN=8'h87;
            BLU=8'h63;
        end
        2504:
        begin
            RED=8'h7C;
            GRN=8'h81;
            BLU=8'h5B;
        end
        2505:
        begin
            RED=8'hB8;
            GRN=8'hA2;
            BLU=8'h73;
        end
        2506:
        begin
            RED=8'hDF;
            GRN=8'hBD;
            BLU=8'h8A;
        end
        2507:
        begin
            RED=8'hD1;
            GRN=8'hA6;
            BLU=8'h74;
        end
        2508:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h88;
        end
        2509:
        begin
            RED=8'hEE;
            GRN=8'hC1;
            BLU=8'h84;
        end
        2510:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h83;
        end
        2511:
        begin
            RED=8'hE3;
            GRN=8'hBB;
            BLU=8'h7D;
        end
        2512:
        begin
            RED=8'hC6;
            GRN=8'h9D;
            BLU=8'h61;
        end
        2513:
        begin
            RED=8'hDB;
            GRN=8'hB1;
            BLU=8'h77;
        end
        2514:
        begin
            RED=8'hEB;
            GRN=8'hBD;
            BLU=8'h85;
        end
        2515:
        begin
            RED=8'hEE;
            GRN=8'hBE;
            BLU=8'h85;
        end
        2516:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h83;
        end
        2517:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h80;
        end
        2518:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h7E;
        end
        2519:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        2520:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        2521:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h82;
        end
        2522:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h81;
        end
        2523:
        begin
            RED=8'hE7;
            GRN=8'hBA;
            BLU=8'h7F;
        end
        2524:
        begin
            RED=8'hC9;
            GRN=8'h9E;
            BLU=8'h6B;
        end
        2525:
        begin
            RED=8'hEB;
            GRN=8'hC0;
            BLU=8'h8A;
        end
        2526:
        begin
            RED=8'hEB;
            GRN=8'hC2;
            BLU=8'h83;
        end
        2527:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h7A;
        end
        2528:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        2529:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        2530:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        2531:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        2532:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        2533:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2534:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2535:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2536:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2537:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        2538:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2539:
        begin
            RED=8'hEC;
            GRN=8'hBE;
            BLU=8'h82;
        end
        2540:
        begin
            RED=8'hEF;
            GRN=8'hC1;
            BLU=8'h87;
        end
        2541:
        begin
            RED=8'hDF;
            GRN=8'hAF;
            BLU=8'h7B;
        end
        2542:
        begin
            RED=8'hE0;
            GRN=8'hB5;
            BLU=8'h82;
        end
        2543:
        begin
            RED=8'hD6;
            GRN=8'hBB;
            BLU=8'h87;
        end
        2544:
        begin
            RED=8'h81;
            GRN=8'h77;
            BLU=8'h5E;
        end
        2545:
        begin
            RED=8'h7D;
            GRN=8'h83;
            BLU=8'h69;
        end
        2546:
        begin
            RED=8'h7C;
            GRN=8'h84;
            BLU=8'h63;
        end
        2547:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2548:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2549:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2550:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2551:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        2552:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h63;
        end
        2553:
        begin
            RED=8'h7B;
            GRN=8'h84;
            BLU=8'h69;
        end
        2554:
        begin
            RED=8'h54;
            GRN=8'h5D;
            BLU=8'h4C;
        end
        2555:
        begin
            RED=8'h2F;
            GRN=8'h33;
            BLU=8'h29;
        end
        2556:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2557:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2558:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2559:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2560:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2561:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2562:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2563:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2564:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h64;
        end
        2565:
        begin
            RED=8'h7C;
            GRN=8'h84;
            BLU=8'h65;
        end
        2566:
        begin
            RED=8'h82;
            GRN=8'h81;
            BLU=8'h63;
        end
        2567:
        begin
            RED=8'h79;
            GRN=8'h87;
            BLU=8'h63;
        end
        2568:
        begin
            RED=8'h7C;
            GRN=8'h89;
            BLU=8'h66;
        end
        2569:
        begin
            RED=8'h7E;
            GRN=8'h74;
            BLU=8'h52;
        end
        2570:
        begin
            RED=8'hB5;
            GRN=8'h98;
            BLU=8'h74;
        end
        2571:
        begin
            RED=8'hC4;
            GRN=8'h9C;
            BLU=8'h6E;
        end
        2572:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h88;
        end
        2573:
        begin
            RED=8'hEA;
            GRN=8'hC2;
            BLU=8'h86;
        end
        2574:
        begin
            RED=8'hDB;
            GRN=8'hB2;
            BLU=8'h7F;
        end
        2575:
        begin
            RED=8'hCB;
            GRN=8'hA2;
            BLU=8'h6C;
        end
        2576:
        begin
            RED=8'hE9;
            GRN=8'hC1;
            BLU=8'h85;
        end
        2577:
        begin
            RED=8'hE9;
            GRN=8'hC2;
            BLU=8'h80;
        end
        2578:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h7F;
        end
        2579:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h7F;
        end
        2580:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        2581:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h83;
        end
        2582:
        begin
            RED=8'hEA;
            GRN=8'hC0;
            BLU=8'h83;
        end
        2583:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        2584:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h82;
        end
        2585:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h83;
        end
        2586:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        2587:
        begin
            RED=8'hEA;
            GRN=8'hBE;
            BLU=8'h7D;
        end
        2588:
        begin
            RED=8'hE6;
            GRN=8'hBB;
            BLU=8'h84;
        end
        2589:
        begin
            RED=8'hC9;
            GRN=8'h9D;
            BLU=8'h6B;
        end
        2590:
        begin
            RED=8'hE9;
            GRN=8'hBE;
            BLU=8'h86;
        end
        2591:
        begin
            RED=8'hEC;
            GRN=8'hC3;
            BLU=8'h80;
        end
        2592:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        2593:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        2594:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        2595:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        2596:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        2597:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2598:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2599:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2600:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2601:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        2602:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2603:
        begin
            RED=8'hED;
            GRN=8'hBE;
            BLU=8'h84;
        end
        2604:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h8A;
        end
        2605:
        begin
            RED=8'hD8;
            GRN=8'hAA;
            BLU=8'h75;
        end
        2606:
        begin
            RED=8'hE1;
            GRN=8'hBD;
            BLU=8'h8A;
        end
        2607:
        begin
            RED=8'h95;
            GRN=8'h84;
            BLU=8'h65;
        end
        2608:
        begin
            RED=8'h80;
            GRN=8'h82;
            BLU=8'h5C;
        end
        2609:
        begin
            RED=8'h80;
            GRN=8'h86;
            BLU=8'h65;
        end
        2610:
        begin
            RED=8'h7D;
            GRN=8'h82;
            BLU=8'h64;
        end
        2611:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2612:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2613:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2614:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2615:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        2616:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h63;
        end
        2617:
        begin
            RED=8'h7B;
            GRN=8'h84;
            BLU=8'h69;
        end
        2618:
        begin
            RED=8'h54;
            GRN=8'h5D;
            BLU=8'h4C;
        end
        2619:
        begin
            RED=8'h2F;
            GRN=8'h33;
            BLU=8'h29;
        end
        2620:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2621:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2622:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2623:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2624:
        begin
            RED=8'h7E;
            GRN=8'h84;
            BLU=8'h62;
        end
        2625:
        begin
            RED=8'h7E;
            GRN=8'h84;
            BLU=8'h62;
        end
        2626:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2627:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        2628:
        begin
            RED=8'h7F;
            GRN=8'h82;
            BLU=8'h65;
        end
        2629:
        begin
            RED=8'h82;
            GRN=8'h81;
            BLU=8'h66;
        end
        2630:
        begin
            RED=8'h81;
            GRN=8'h82;
            BLU=8'h62;
        end
        2631:
        begin
            RED=8'h7E;
            GRN=8'h84;
            BLU=8'h62;
        end
        2632:
        begin
            RED=8'h7E;
            GRN=8'h81;
            BLU=8'h62;
        end
        2633:
        begin
            RED=8'h8C;
            GRN=8'h77;
            BLU=8'h53;
        end
        2634:
        begin
            RED=8'hE3;
            GRN=8'hBD;
            BLU=8'h8D;
        end
        2635:
        begin
            RED=8'hDF;
            GRN=8'hB5;
            BLU=8'h7A;
        end
        2636:
        begin
            RED=8'hC2;
            GRN=8'h99;
            BLU=8'h61;
        end
        2637:
        begin
            RED=8'hC1;
            GRN=8'h9B;
            BLU=8'h68;
        end
        2638:
        begin
            RED=8'hD9;
            GRN=8'hAC;
            BLU=8'h75;
        end
        2639:
        begin
            RED=8'hEE;
            GRN=8'hC1;
            BLU=8'h87;
        end
        2640:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h84;
        end
        2641:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h83;
        end
        2642:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h80;
        end
        2643:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2644:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2645:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2646:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2647:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2648:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h80;
        end
        2649:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h80;
        end
        2650:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        2651:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2652:
        begin
            RED=8'hEF;
            GRN=8'hC2;
            BLU=8'h83;
        end
        2653:
        begin
            RED=8'hE6;
            GRN=8'hB9;
            BLU=8'h7C;
        end
        2654:
        begin
            RED=8'hD0;
            GRN=8'hA4;
            BLU=8'h65;
        end
        2655:
        begin
            RED=8'hEA;
            GRN=8'hBE;
            BLU=8'h7D;
        end
        2656:
        begin
            RED=8'hEE;
            GRN=8'hC1;
            BLU=8'h7F;
        end
        2657:
        begin
            RED=8'hEE;
            GRN=8'hC1;
            BLU=8'h7E;
        end
        2658:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h7D;
        end
        2659:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        2660:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        2661:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2662:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2663:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2664:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2665:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2666:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h7E;
        end
        2667:
        begin
            RED=8'hEC;
            GRN=8'hC1;
            BLU=8'h7E;
        end
        2668:
        begin
            RED=8'hEA;
            GRN=8'hC0;
            BLU=8'h88;
        end
        2669:
        begin
            RED=8'hC6;
            GRN=8'h9B;
            BLU=8'h68;
        end
        2670:
        begin
            RED=8'hDB;
            GRN=8'hBD;
            BLU=8'h88;
        end
        2671:
        begin
            RED=8'h7C;
            GRN=8'h7A;
            BLU=8'h5E;
        end
        2672:
        begin
            RED=8'h80;
            GRN=8'h83;
            BLU=8'h63;
        end
        2673:
        begin
            RED=8'h81;
            GRN=8'h82;
            BLU=8'h63;
        end
        2674:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h64;
        end
        2675:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2676:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2677:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2678:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2679:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h65;
        end
        2680:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h64;
        end
        2681:
        begin
            RED=8'h7C;
            GRN=8'h84;
            BLU=8'h6A;
        end
        2682:
        begin
            RED=8'h57;
            GRN=8'h5E;
            BLU=8'h4F;
        end
        2683:
        begin
            RED=8'h2E;
            GRN=8'h32;
            BLU=8'h29;
        end
        2684:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2685:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2686:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2687:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2688:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        2689:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2690:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2691:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2692:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h63;
        end
        2693:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h62;
        end
        2694:
        begin
            RED=8'h7C;
            GRN=8'h84;
            BLU=8'h63;
        end
        2695:
        begin
            RED=8'h7D;
            GRN=8'h82;
            BLU=8'h63;
        end
        2696:
        begin
            RED=8'h80;
            GRN=8'h7F;
            BLU=8'h63;
        end
        2697:
        begin
            RED=8'hBA;
            GRN=8'hA0;
            BLU=8'h72;
        end
        2698:
        begin
            RED=8'hE9;
            GRN=8'hC1;
            BLU=8'h84;
        end
        2699:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        2700:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h82;
        end
        2701:
        begin
            RED=8'hE8;
            GRN=8'hC0;
            BLU=8'h89;
        end
        2702:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h85;
        end
        2703:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h85;
        end
        2704:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h83;
        end
        2705:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h83;
        end
        2706:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        2707:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2708:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2709:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2710:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2711:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2712:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2713:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2714:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2715:
        begin
            RED=8'hEE;
            GRN=8'hC1;
            BLU=8'h80;
        end
        2716:
        begin
            RED=8'hEE;
            GRN=8'hC1;
            BLU=8'h80;
        end
        2717:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2718:
        begin
            RED=8'hEB;
            GRN=8'hBE;
            BLU=8'h7D;
        end
        2719:
        begin
            RED=8'hD9;
            GRN=8'hAC;
            BLU=8'h6C;
        end
        2720:
        begin
            RED=8'hDD;
            GRN=8'hB0;
            BLU=8'h74;
        end
        2721:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h82;
        end
        2722:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h7F;
        end
        2723:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7C;
        end
        2724:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7C;
        end
        2725:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2726:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2727:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2728:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2729:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h81;
        end
        2730:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h7F;
        end
        2731:
        begin
            RED=8'hE5;
            GRN=8'hBB;
            BLU=8'h7A;
        end
        2732:
        begin
            RED=8'hDE;
            GRN=8'hB5;
            BLU=8'h7C;
        end
        2733:
        begin
            RED=8'hC9;
            GRN=8'hA0;
            BLU=8'h6C;
        end
        2734:
        begin
            RED=8'hBF;
            GRN=8'hA5;
            BLU=8'h76;
        end
        2735:
        begin
            RED=8'h7C;
            GRN=8'h7E;
            BLU=8'h63;
        end
        2736:
        begin
            RED=8'h80;
            GRN=8'h82;
            BLU=8'h65;
        end
        2737:
        begin
            RED=8'h80;
            GRN=8'h82;
            BLU=8'h63;
        end
        2738:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        2739:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2740:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2741:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2742:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2743:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        2744:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h63;
        end
        2745:
        begin
            RED=8'h7C;
            GRN=8'h85;
            BLU=8'h69;
        end
        2746:
        begin
            RED=8'h57;
            GRN=8'h5F;
            BLU=8'h4E;
        end
        2747:
        begin
            RED=8'h2E;
            GRN=8'h32;
            BLU=8'h28;
        end
        2748:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2749:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2750:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2751:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2752:
        begin
            RED=8'h7D;
            GRN=8'h81;
            BLU=8'h69;
        end
        2753:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h68;
        end
        2754:
        begin
            RED=8'h7D;
            GRN=8'h82;
            BLU=8'h65;
        end
        2755:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2756:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h61;
        end
        2757:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h5F;
        end
        2758:
        begin
            RED=8'h79;
            GRN=8'h86;
            BLU=8'h64;
        end
        2759:
        begin
            RED=8'h7D;
            GRN=8'h83;
            BLU=8'h64;
        end
        2760:
        begin
            RED=8'h82;
            GRN=8'h77;
            BLU=8'h58;
        end
        2761:
        begin
            RED=8'hD9;
            GRN=8'hBA;
            BLU=8'h84;
        end
        2762:
        begin
            RED=8'hED;
            GRN=8'hC3;
            BLU=8'h7F;
        end
        2763:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7A;
        end
        2764:
        begin
            RED=8'hEB;
            GRN=8'hC0;
            BLU=8'h7C;
        end
        2765:
        begin
            RED=8'hE9;
            GRN=8'hC2;
            BLU=8'h81;
        end
        2766:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h82;
        end
        2767:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h83;
        end
        2768:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h83;
        end
        2769:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h82;
        end
        2770:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2771:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2772:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2773:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2774:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2775:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2776:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2777:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2778:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2779:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2780:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2781:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2782:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        2783:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2784:
        begin
            RED=8'hE3;
            GRN=8'hB5;
            BLU=8'h7C;
        end
        2785:
        begin
            RED=8'hD1;
            GRN=8'hA5;
            BLU=8'h6A;
        end
        2786:
        begin
            RED=8'hEB;
            GRN=8'hBD;
            BLU=8'h7F;
        end
        2787:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        2788:
        begin
            RED=8'hEE;
            GRN=8'hC1;
            BLU=8'h7E;
        end
        2789:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2790:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2791:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2792:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2793:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h82;
        end
        2794:
        begin
            RED=8'hEC;
            GRN=8'hBE;
            BLU=8'h83;
        end
        2795:
        begin
            RED=8'hD9;
            GRN=8'hAE;
            BLU=8'h74;
        end
        2796:
        begin
            RED=8'hD6;
            GRN=8'hAD;
            BLU=8'h75;
        end
        2797:
        begin
            RED=8'hE6;
            GRN=8'hC0;
            BLU=8'h8B;
        end
        2798:
        begin
            RED=8'h9B;
            GRN=8'h8A;
            BLU=8'h64;
        end
        2799:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h6A;
        end
        2800:
        begin
            RED=8'h7F;
            GRN=8'h82;
            BLU=8'h65;
        end
        2801:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2802:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h64;
        end
        2803:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2804:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2805:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2806:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2807:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2808:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h62;
        end
        2809:
        begin
            RED=8'h7C;
            GRN=8'h85;
            BLU=8'h68;
        end
        2810:
        begin
            RED=8'h57;
            GRN=8'h60;
            BLU=8'h4D;
        end
        2811:
        begin
            RED=8'h2E;
            GRN=8'h32;
            BLU=8'h28;
        end
        2812:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2813:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2814:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2815:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2816:
        begin
            RED=8'h7E;
            GRN=8'h81;
            BLU=8'h6F;
        end
        2817:
        begin
            RED=8'h80;
            GRN=8'h83;
            BLU=8'h6D;
        end
        2818:
        begin
            RED=8'h7D;
            GRN=8'h81;
            BLU=8'h67;
        end
        2819:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2820:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h62;
        end
        2821:
        begin
            RED=8'h80;
            GRN=8'h82;
            BLU=8'h66;
        end
        2822:
        begin
            RED=8'h7B;
            GRN=8'h84;
            BLU=8'h69;
        end
        2823:
        begin
            RED=8'h7F;
            GRN=8'h7F;
            BLU=8'h60;
        end
        2824:
        begin
            RED=8'hA3;
            GRN=8'h8B;
            BLU=8'h61;
        end
        2825:
        begin
            RED=8'hE7;
            GRN=8'hC1;
            BLU=8'h84;
        end
        2826:
        begin
            RED=8'hEC;
            GRN=8'hC1;
            BLU=8'h7D;
        end
        2827:
        begin
            RED=8'hF0;
            GRN=8'hBF;
            BLU=8'h7D;
        end
        2828:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        2829:
        begin
            RED=8'hEA;
            GRN=8'hC2;
            BLU=8'h7D;
        end
        2830:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2831:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2832:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2833:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2834:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2835:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2836:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2837:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2838:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2839:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2840:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2841:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2842:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2843:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2844:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2845:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2846:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2847:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2848:
        begin
            RED=8'hEF;
            GRN=8'hC1;
            BLU=8'h82;
        end
        2849:
        begin
            RED=8'hEB;
            GRN=8'hBE;
            BLU=8'h80;
        end
        2850:
        begin
            RED=8'hD4;
            GRN=8'hA6;
            BLU=8'h6B;
        end
        2851:
        begin
            RED=8'hE2;
            GRN=8'hB3;
            BLU=8'h79;
        end
        2852:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h84;
        end
        2853:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2854:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2855:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2856:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2857:
        begin
            RED=8'hEC;
            GRN=8'hBE;
            BLU=8'h82;
        end
        2858:
        begin
            RED=8'hD7;
            GRN=8'hA9;
            BLU=8'h74;
        end
        2859:
        begin
            RED=8'hEB;
            GRN=8'hBF;
            BLU=8'h8C;
        end
        2860:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h89;
        end
        2861:
        begin
            RED=8'hE1;
            GRN=8'hBE;
            BLU=8'h87;
        end
        2862:
        begin
            RED=8'h81;
            GRN=8'h77;
            BLU=8'h5C;
        end
        2863:
        begin
            RED=8'h7D;
            GRN=8'h83;
            BLU=8'h6E;
        end
        2864:
        begin
            RED=8'h7F;
            GRN=8'h82;
            BLU=8'h63;
        end
        2865:
        begin
            RED=8'h7C;
            GRN=8'h85;
            BLU=8'h63;
        end
        2866:
        begin
            RED=8'h7C;
            GRN=8'h84;
            BLU=8'h64;
        end
        2867:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2868:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2869:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2870:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2871:
        begin
            RED=8'h7E;
            GRN=8'h84;
            BLU=8'h61;
        end
        2872:
        begin
            RED=8'h7D;
            GRN=8'h85;
            BLU=8'h60;
        end
        2873:
        begin
            RED=8'h7C;
            GRN=8'h85;
            BLU=8'h66;
        end
        2874:
        begin
            RED=8'h57;
            GRN=8'h60;
            BLU=8'h4B;
        end
        2875:
        begin
            RED=8'h2E;
            GRN=8'h32;
            BLU=8'h27;
        end
        2876:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2877:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2878:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2879:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2880:
        begin
            RED=8'h3F;
            GRN=8'h42;
            BLU=8'h34;
        end
        2881:
        begin
            RED=8'h6D;
            GRN=8'h70;
            BLU=8'h60;
        end
        2882:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h6C;
        end
        2883:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h65;
        end
        2884:
        begin
            RED=8'h80;
            GRN=8'h83;
            BLU=8'h63;
        end
        2885:
        begin
            RED=8'h81;
            GRN=8'h80;
            BLU=8'h6A;
        end
        2886:
        begin
            RED=8'h7D;
            GRN=8'h7E;
            BLU=8'h66;
        end
        2887:
        begin
            RED=8'h83;
            GRN=8'h75;
            BLU=8'h52;
        end
        2888:
        begin
            RED=8'hE2;
            GRN=8'hBA;
            BLU=8'h85;
        end
        2889:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2890:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2891:
        begin
            RED=8'hF0;
            GRN=8'hBE;
            BLU=8'h81;
        end
        2892:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h80;
        end
        2893:
        begin
            RED=8'hEC;
            GRN=8'hC1;
            BLU=8'h7F;
        end
        2894:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h82;
        end
        2895:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2896:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h7F;
        end
        2897:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h7F;
        end
        2898:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h80;
        end
        2899:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2900:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2901:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2902:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2903:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2904:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2905:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2906:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        2907:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2908:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        2909:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        2910:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2911:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2912:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7C;
        end
        2913:
        begin
            RED=8'hEB;
            GRN=8'hBE;
            BLU=8'h7C;
        end
        2914:
        begin
            RED=8'hEC;
            GRN=8'hBE;
            BLU=8'h84;
        end
        2915:
        begin
            RED=8'hD6;
            GRN=8'hA7;
            BLU=8'h72;
        end
        2916:
        begin
            RED=8'hE1;
            GRN=8'hB2;
            BLU=8'h7C;
        end
        2917:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2918:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2919:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2920:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2921:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h81;
        end
        2922:
        begin
            RED=8'hC6;
            GRN=8'h98;
            BLU=8'h65;
        end
        2923:
        begin
            RED=8'hE4;
            GRN=8'hB8;
            BLU=8'h87;
        end
        2924:
        begin
            RED=8'hE3;
            GRN=8'hBE;
            BLU=8'h8A;
        end
        2925:
        begin
            RED=8'hA3;
            GRN=8'h8B;
            BLU=8'h59;
        end
        2926:
        begin
            RED=8'h83;
            GRN=8'h80;
            BLU=8'h67;
        end
        2927:
        begin
            RED=8'h7D;
            GRN=8'h85;
            BLU=8'h6E;
        end
        2928:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2929:
        begin
            RED=8'h7B;
            GRN=8'h84;
            BLU=8'h63;
        end
        2930:
        begin
            RED=8'h7C;
            GRN=8'h84;
            BLU=8'h65;
        end
        2931:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2932:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2933:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2934:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2935:
        begin
            RED=8'h7E;
            GRN=8'h84;
            BLU=8'h60;
        end
        2936:
        begin
            RED=8'h7D;
            GRN=8'h85;
            BLU=8'h5E;
        end
        2937:
        begin
            RED=8'h7C;
            GRN=8'h85;
            BLU=8'h65;
        end
        2938:
        begin
            RED=8'h57;
            GRN=8'h60;
            BLU=8'h4A;
        end
        2939:
        begin
            RED=8'h2E;
            GRN=8'h32;
            BLU=8'h26;
        end
        2940:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2941:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2942:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2943:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        2944:
        begin
            RED=8'h2D;
            GRN=8'h33;
            BLU=8'h29;
        end
        2945:
        begin
            RED=8'h2C;
            GRN=8'h2F;
            BLU=8'h28;
        end
        2946:
        begin
            RED=8'h47;
            GRN=8'h49;
            BLU=8'h3D;
        end
        2947:
        begin
            RED=8'h76;
            GRN=8'h78;
            BLU=8'h61;
        end
        2948:
        begin
            RED=8'h7E;
            GRN=8'h7D;
            BLU=8'h5B;
        end
        2949:
        begin
            RED=8'h91;
            GRN=8'h86;
            BLU=8'h5A;
        end
        2950:
        begin
            RED=8'hAE;
            GRN=8'h9A;
            BLU=8'h68;
        end
        2951:
        begin
            RED=8'hE1;
            GRN=8'hBE;
            BLU=8'h85;
        end
        2952:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h7F;
        end
        2953:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h7F;
        end
        2954:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h82;
        end
        2955:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h82;
        end
        2956:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h82;
        end
        2957:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h82;
        end
        2958:
        begin
            RED=8'hE9;
            GRN=8'hC1;
            BLU=8'h84;
        end
        2959:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h81;
        end
        2960:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        2961:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        2962:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2963:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2964:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2965:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2966:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2967:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2968:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2969:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2970:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2971:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h7E;
        end
        2972:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h7D;
        end
        2973:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h7E;
        end
        2974:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2975:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2976:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2977:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2978:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2979:
        begin
            RED=8'hEF;
            GRN=8'hC2;
            BLU=8'h82;
        end
        2980:
        begin
            RED=8'hD5;
            GRN=8'hA9;
            BLU=8'h68;
        end
        2981:
        begin
            RED=8'hE4;
            GRN=8'hB8;
            BLU=8'h77;
        end
        2982:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2983:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2984:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        2985:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h7A;
        end
        2986:
        begin
            RED=8'hEA;
            GRN=8'hBF;
            BLU=8'h85;
        end
        2987:
        begin
            RED=8'hD1;
            GRN=8'hA6;
            BLU=8'h72;
        end
        2988:
        begin
            RED=8'hA2;
            GRN=8'h89;
            BLU=8'h62;
        end
        2989:
        begin
            RED=8'h73;
            GRN=8'h78;
            BLU=8'h60;
        end
        2990:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h64;
        end
        2991:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h66;
        end
        2992:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h67;
        end
        2993:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h67;
        end
        2994:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h65;
        end
        2995:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2996:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2997:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2998:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        2999:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h62;
        end
        3000:
        begin
            RED=8'h7D;
            GRN=8'h85;
            BLU=8'h60;
        end
        3001:
        begin
            RED=8'h7C;
            GRN=8'h86;
            BLU=8'h65;
        end
        3002:
        begin
            RED=8'h58;
            GRN=8'h62;
            BLU=8'h49;
        end
        3003:
        begin
            RED=8'h2D;
            GRN=8'h32;
            BLU=8'h25;
        end
        3004:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3005:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3006:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3007:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3008:
        begin
            RED=8'h2E;
            GRN=8'h33;
            BLU=8'h28;
        end
        3009:
        begin
            RED=8'h2E;
            GRN=8'h31;
            BLU=8'h29;
        end
        3010:
        begin
            RED=8'h2D;
            GRN=8'h2F;
            BLU=8'h26;
        end
        3011:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h1F;
        end
        3012:
        begin
            RED=8'hAA;
            GRN=8'hA2;
            BLU=8'h7E;
        end
        3013:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h7D;
        end
        3014:
        begin
            RED=8'hEC;
            GRN=8'hC2;
            BLU=8'h7F;
        end
        3015:
        begin
            RED=8'hEA;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        3016:
        begin
            RED=8'hE9;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3017:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3018:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        3019:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        3020:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        3021:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h7C;
        end
        3022:
        begin
            RED=8'hF0;
            GRN=8'hC0;
            BLU=8'h76;
        end
        3023:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h7B;
        end
        3024:
        begin
            RED=8'hEA;
            GRN=8'hC2;
            BLU=8'h7D;
        end
        3025:
        begin
            RED=8'hE9;
            GRN=8'hC2;
            BLU=8'h7E;
        end
        3026:
        begin
            RED=8'hEB;
            GRN=8'hC1;
            BLU=8'h7C;
        end
        3027:
        begin
            RED=8'hEC;
            GRN=8'hC1;
            BLU=8'h7C;
        end
        3028:
        begin
            RED=8'hEC;
            GRN=8'hC1;
            BLU=8'h7C;
        end
        3029:
        begin
            RED=8'hEC;
            GRN=8'hC1;
            BLU=8'h7C;
        end
        3030:
        begin
            RED=8'hEC;
            GRN=8'hC1;
            BLU=8'h7C;
        end
        3031:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7C;
        end
        3032:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7C;
        end
        3033:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7C;
        end
        3034:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7C;
        end
        3035:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h81;
        end
        3036:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h87;
        end
        3037:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h84;
        end
        3038:
        begin
            RED=8'hEB;
            GRN=8'hC1;
            BLU=8'h81;
        end
        3039:
        begin
            RED=8'hEB;
            GRN=8'hC1;
            BLU=8'h80;
        end
        3040:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3041:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3042:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3043:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3044:
        begin
            RED=8'hEB;
            GRN=8'hBE;
            BLU=8'h7D;
        end
        3045:
        begin
            RED=8'hD1;
            GRN=8'hA4;
            BLU=8'h63;
        end
        3046:
        begin
            RED=8'hEF;
            GRN=8'hC2;
            BLU=8'h81;
        end
        3047:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3048:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3049:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h77;
        end
        3050:
        begin
            RED=8'hEC;
            GRN=8'hC4;
            BLU=8'h82;
        end
        3051:
        begin
            RED=8'hEB;
            GRN=8'hBF;
            BLU=8'h86;
        end
        3052:
        begin
            RED=8'hCC;
            GRN=8'hB0;
            BLU=8'h8A;
        end
        3053:
        begin
            RED=8'hDC;
            GRN=8'hDC;
            BLU=8'hD0;
        end
        3054:
        begin
            RED=8'h90;
            GRN=8'h92;
            BLU=8'h86;
        end
        3055:
        begin
            RED=8'h78;
            GRN=8'h7B;
            BLU=8'h6A;
        end
        3056:
        begin
            RED=8'h7E;
            GRN=8'h81;
            BLU=8'h6A;
        end
        3057:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h65;
        end
        3058:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        3059:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        3060:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        3061:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        3062:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        3063:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h62;
        end
        3064:
        begin
            RED=8'h7D;
            GRN=8'h85;
            BLU=8'h60;
        end
        3065:
        begin
            RED=8'h7C;
            GRN=8'h86;
            BLU=8'h65;
        end
        3066:
        begin
            RED=8'h58;
            GRN=8'h62;
            BLU=8'h49;
        end
        3067:
        begin
            RED=8'h2D;
            GRN=8'h32;
            BLU=8'h25;
        end
        3068:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3069:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3070:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3071:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3072:
        begin
            RED=8'h2D;
            GRN=8'h33;
            BLU=8'h26;
        end
        3073:
        begin
            RED=8'h2F;
            GRN=8'h32;
            BLU=8'h2A;
        end
        3074:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h29;
        end
        3075:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h22;
        end
        3076:
        begin
            RED=8'h44;
            GRN=8'h3F;
            BLU=8'h27;
        end
        3077:
        begin
            RED=8'hAA;
            GRN=8'h93;
            BLU=8'h68;
        end
        3078:
        begin
            RED=8'hDA;
            GRN=8'hBC;
            BLU=8'h8A;
        end
        3079:
        begin
            RED=8'hE9;
            GRN=8'hC1;
            BLU=8'h85;
        end
        3080:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h7B;
        end
        3081:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h7C;
        end
        3082:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        3083:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        3084:
        begin
            RED=8'hEF;
            GRN=8'hC1;
            BLU=8'h7E;
        end
        3085:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h7C;
        end
        3086:
        begin
            RED=8'hEF;
            GRN=8'hBD;
            BLU=8'h7D;
        end
        3087:
        begin
            RED=8'hE9;
            GRN=8'hC1;
            BLU=8'h89;
        end
        3088:
        begin
            RED=8'hE3;
            GRN=8'hBF;
            BLU=8'h8B;
        end
        3089:
        begin
            RED=8'hDB;
            GRN=8'hB4;
            BLU=8'h7C;
        end
        3090:
        begin
            RED=8'hDB;
            GRN=8'hB1;
            BLU=8'h78;
        end
        3091:
        begin
            RED=8'hDB;
            GRN=8'hB1;
            BLU=8'h78;
        end
        3092:
        begin
            RED=8'hE0;
            GRN=8'hB6;
            BLU=8'h7C;
        end
        3093:
        begin
            RED=8'hE4;
            GRN=8'hBA;
            BLU=8'h81;
        end
        3094:
        begin
            RED=8'hE0;
            GRN=8'hB6;
            BLU=8'h7C;
        end
        3095:
        begin
            RED=8'hDA;
            GRN=8'hAC;
            BLU=8'h74;
        end
        3096:
        begin
            RED=8'hD3;
            GRN=8'hA4;
            BLU=8'h6C;
        end
        3097:
        begin
            RED=8'hD6;
            GRN=8'hA7;
            BLU=8'h70;
        end
        3098:
        begin
            RED=8'hD0;
            GRN=8'hA1;
            BLU=8'h6A;
        end
        3099:
        begin
            RED=8'hCD;
            GRN=8'h9D;
            BLU=8'h67;
        end
        3100:
        begin
            RED=8'hD2;
            GRN=8'hA3;
            BLU=8'h6E;
        end
        3101:
        begin
            RED=8'hDD;
            GRN=8'hB1;
            BLU=8'h7B;
        end
        3102:
        begin
            RED=8'hDF;
            GRN=8'hB7;
            BLU=8'h7F;
        end
        3103:
        begin
            RED=8'hE2;
            GRN=8'hBB;
            BLU=8'h83;
        end
        3104:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h81;
        end
        3105:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3106:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3107:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3108:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3109:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        3110:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3111:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3112:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3113:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h7C;
        end
        3114:
        begin
            RED=8'hEA;
            GRN=8'hC2;
            BLU=8'h7F;
        end
        3115:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h82;
        end
        3116:
        begin
            RED=8'hD9;
            GRN=8'hB8;
            BLU=8'h8F;
        end
        3117:
        begin
            RED=8'hEF;
            GRN=8'hEC;
            BLU=8'hE3;
        end
        3118:
        begin
            RED=8'hF6;
            GRN=8'hF6;
            BLU=8'hF7;
        end
        3119:
        begin
            RED=8'hCB;
            GRN=8'hCC;
            BLU=8'hC5;
        end
        3120:
        begin
            RED=8'h79;
            GRN=8'h7C;
            BLU=8'h6C;
        end
        3121:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h6B;
        end
        3122:
        begin
            RED=8'h7D;
            GRN=8'h82;
            BLU=8'h64;
        end
        3123:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        3124:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        3125:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        3126:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        3127:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h62;
        end
        3128:
        begin
            RED=8'h7D;
            GRN=8'h85;
            BLU=8'h60;
        end
        3129:
        begin
            RED=8'h7C;
            GRN=8'h85;
            BLU=8'h64;
        end
        3130:
        begin
            RED=8'h58;
            GRN=8'h62;
            BLU=8'h49;
        end
        3131:
        begin
            RED=8'h2E;
            GRN=8'h32;
            BLU=8'h25;
        end
        3132:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3133:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3134:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3135:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3136:
        begin
            RED=8'h2D;
            GRN=8'h33;
            BLU=8'h25;
        end
        3137:
        begin
            RED=8'h2F;
            GRN=8'h32;
            BLU=8'h2A;
        end
        3138:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h2B;
        end
        3139:
        begin
            RED=8'h30;
            GRN=8'h30;
            BLU=8'h27;
        end
        3140:
        begin
            RED=8'h2E;
            GRN=8'h2D;
            BLU=8'h1F;
        end
        3141:
        begin
            RED=8'h33;
            GRN=8'h31;
            BLU=8'h22;
        end
        3142:
        begin
            RED=8'h46;
            GRN=8'h3E;
            BLU=8'h29;
        end
        3143:
        begin
            RED=8'h73;
            GRN=8'h66;
            BLU=8'h48;
        end
        3144:
        begin
            RED=8'hA7;
            GRN=8'h94;
            BLU=8'h6D;
        end
        3145:
        begin
            RED=8'hC1;
            GRN=8'hAD;
            BLU=8'h7E;
        end
        3146:
        begin
            RED=8'hC2;
            GRN=8'hAD;
            BLU=8'h7D;
        end
        3147:
        begin
            RED=8'hBF;
            GRN=8'hAB;
            BLU=8'h7A;
        end
        3148:
        begin
            RED=8'hB8;
            GRN=8'hA4;
            BLU=8'h73;
        end
        3149:
        begin
            RED=8'hAD;
            GRN=8'h99;
            BLU=8'h69;
        end
        3150:
        begin
            RED=8'h93;
            GRN=8'h82;
            BLU=8'h57;
        end
        3151:
        begin
            RED=8'h86;
            GRN=8'h7F;
            BLU=8'h5B;
        end
        3152:
        begin
            RED=8'h7E;
            GRN=8'h78;
            BLU=8'h56;
        end
        3153:
        begin
            RED=8'h87;
            GRN=8'h75;
            BLU=8'h4C;
        end
        3154:
        begin
            RED=8'hDC;
            GRN=8'hBA;
            BLU=8'h83;
        end
        3155:
        begin
            RED=8'hDF;
            GRN=8'hB7;
            BLU=8'h7A;
        end
        3156:
        begin
            RED=8'hDB;
            GRN=8'hB2;
            BLU=8'h76;
        end
        3157:
        begin
            RED=8'hD5;
            GRN=8'hAD;
            BLU=8'h71;
        end
        3158:
        begin
            RED=8'hDB;
            GRN=8'hB2;
            BLU=8'h76;
        end
        3159:
        begin
            RED=8'hE6;
            GRN=8'hB8;
            BLU=8'h7D;
        end
        3160:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h85;
        end
        3161:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h84;
        end
        3162:
        begin
            RED=8'hEF;
            GRN=8'hC1;
            BLU=8'h86;
        end
        3163:
        begin
            RED=8'hF0;
            GRN=8'hC1;
            BLU=8'h86;
        end
        3164:
        begin
            RED=8'hEA;
            GRN=8'hBB;
            BLU=8'h82;
        end
        3165:
        begin
            RED=8'hDE;
            GRN=8'hB3;
            BLU=8'h7F;
        end
        3166:
        begin
            RED=8'hC0;
            GRN=8'h99;
            BLU=8'h6C;
        end
        3167:
        begin
            RED=8'hB0;
            GRN=8'h8D;
            BLU=8'h62;
        end
        3168:
        begin
            RED=8'hEC;
            GRN=8'hC1;
            BLU=8'h84;
        end
        3169:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3170:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3171:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3172:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3173:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3174:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3175:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3176:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3177:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h84;
        end
        3178:
        begin
            RED=8'hEA;
            GRN=8'hC1;
            BLU=8'h83;
        end
        3179:
        begin
            RED=8'hEF;
            GRN=8'hC0;
            BLU=8'h7C;
        end
        3180:
        begin
            RED=8'hDF;
            GRN=8'hBC;
            BLU=8'h8A;
        end
        3181:
        begin
            RED=8'hDC;
            GRN=8'hD4;
            BLU=8'hC6;
        end
        3182:
        begin
            RED=8'hF9;
            GRN=8'hF8;
            BLU=8'hFC;
        end
        3183:
        begin
            RED=8'hF9;
            GRN=8'hF9;
            BLU=8'hF8;
        end
        3184:
        begin
            RED=8'hE6;
            GRN=8'hE7;
            BLU=8'hE0;
        end
        3185:
        begin
            RED=8'h7E;
            GRN=8'h80;
            BLU=8'h74;
        end
        3186:
        begin
            RED=8'h7B;
            GRN=8'h7F;
            BLU=8'h65;
        end
        3187:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        3188:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        3189:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        3190:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        3191:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h62;
        end
        3192:
        begin
            RED=8'h7D;
            GRN=8'h85;
            BLU=8'h60;
        end
        3193:
        begin
            RED=8'h7C;
            GRN=8'h85;
            BLU=8'h64;
        end
        3194:
        begin
            RED=8'h58;
            GRN=8'h62;
            BLU=8'h49;
        end
        3195:
        begin
            RED=8'h2E;
            GRN=8'h32;
            BLU=8'h25;
        end
        3196:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3197:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3198:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3199:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3200:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h28;
        end
        3201:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3202:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h2B;
        end
        3203:
        begin
            RED=8'h31;
            GRN=8'h31;
            BLU=8'h29;
        end
        3204:
        begin
            RED=8'h30;
            GRN=8'h30;
            BLU=8'h26;
        end
        3205:
        begin
            RED=8'h30;
            GRN=8'h2F;
            BLU=8'h28;
        end
        3206:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h28;
        end
        3207:
        begin
            RED=8'h31;
            GRN=8'h32;
            BLU=8'h26;
        end
        3208:
        begin
            RED=8'h2C;
            GRN=8'h2D;
            BLU=8'h21;
        end
        3209:
        begin
            RED=8'h4A;
            GRN=8'h4C;
            BLU=8'h3A;
        end
        3210:
        begin
            RED=8'h77;
            GRN=8'h78;
            BLU=8'h63;
        end
        3211:
        begin
            RED=8'h7C;
            GRN=8'h7E;
            BLU=8'h65;
        end
        3212:
        begin
            RED=8'h7D;
            GRN=8'h7F;
            BLU=8'h62;
        end
        3213:
        begin
            RED=8'h7F;
            GRN=8'h82;
            BLU=8'h61;
        end
        3214:
        begin
            RED=8'h7E;
            GRN=8'h84;
            BLU=8'h66;
        end
        3215:
        begin
            RED=8'h7C;
            GRN=8'h84;
            BLU=8'h67;
        end
        3216:
        begin
            RED=8'h7F;
            GRN=8'h85;
            BLU=8'h67;
        end
        3217:
        begin
            RED=8'h7B;
            GRN=8'h7C;
            BLU=8'h59;
        end
        3218:
        begin
            RED=8'hCA;
            GRN=8'hB0;
            BLU=8'h7F;
        end
        3219:
        begin
            RED=8'hEC;
            GRN=8'hC1;
            BLU=8'h84;
        end
        3220:
        begin
            RED=8'hEE;
            GRN=8'hC2;
            BLU=8'h81;
        end
        3221:
        begin
            RED=8'hEE;
            GRN=8'hC3;
            BLU=8'h81;
        end
        3222:
        begin
            RED=8'hEB;
            GRN=8'hC2;
            BLU=8'h7F;
        end
        3223:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h7F;
        end
        3224:
        begin
            RED=8'hEE;
            GRN=8'hC1;
            BLU=8'h7F;
        end
        3225:
        begin
            RED=8'hEF;
            GRN=8'hC2;
            BLU=8'h80;
        end
        3226:
        begin
            RED=8'hF0;
            GRN=8'hC3;
            BLU=8'h81;
        end
        3227:
        begin
            RED=8'hEF;
            GRN=8'hC2;
            BLU=8'h80;
        end
        3228:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3229:
        begin
            RED=8'hEB;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        3230:
        begin
            RED=8'hEB;
            GRN=8'hBF;
            BLU=8'h88;
        end
        3231:
        begin
            RED=8'hCD;
            GRN=8'hA1;
            BLU=8'h74;
        end
        3232:
        begin
            RED=8'hE2;
            GRN=8'hB5;
            BLU=8'h78;
        end
        3233:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3234:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3235:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3236:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3237:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h7F;
        end
        3238:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        3239:
        begin
            RED=8'hEB;
            GRN=8'hBF;
            BLU=8'h7C;
        end
        3240:
        begin
            RED=8'hEC;
            GRN=8'hC2;
            BLU=8'h7E;
        end
        3241:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h80;
        end
        3242:
        begin
            RED=8'hE9;
            GRN=8'hC1;
            BLU=8'h85;
        end
        3243:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h80;
        end
        3244:
        begin
            RED=8'hE8;
            GRN=8'hC3;
            BLU=8'h89;
        end
        3245:
        begin
            RED=8'hAF;
            GRN=8'hA2;
            BLU=8'h85;
        end
        3246:
        begin
            RED=8'hED;
            GRN=8'hEF;
            BLU=8'hF3;
        end
        3247:
        begin
            RED=8'hFB;
            GRN=8'hFA;
            BLU=8'hFA;
        end
        3248:
        begin
            RED=8'hFA;
            GRN=8'hF9;
            BLU=8'hF5;
        end
        3249:
        begin
            RED=8'hEE;
            GRN=8'hF0;
            BLU=8'hEC;
        end
        3250:
        begin
            RED=8'h83;
            GRN=8'h87;
            BLU=8'h78;
        end
        3251:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h67;
        end
        3252:
        begin
            RED=8'h7B;
            GRN=8'h81;
            BLU=8'h5F;
        end
        3253:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        3254:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h66;
        end
        3255:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        3256:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h63;
        end
        3257:
        begin
            RED=8'h7C;
            GRN=8'h85;
            BLU=8'h66;
        end
        3258:
        begin
            RED=8'h58;
            GRN=8'h61;
            BLU=8'h4B;
        end
        3259:
        begin
            RED=8'h2D;
            GRN=8'h31;
            BLU=8'h25;
        end
        3260:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h28;
        end
        3261:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3262:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3263:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3264:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3265:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3266:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3267:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3268:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3269:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3270:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3271:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3272:
        begin
            RED=8'h2E;
            GRN=8'h2F;
            BLU=8'h27;
        end
        3273:
        begin
            RED=8'h2C;
            GRN=8'h2F;
            BLU=8'h24;
        end
        3274:
        begin
            RED=8'h31;
            GRN=8'h35;
            BLU=8'h28;
        end
        3275:
        begin
            RED=8'h5D;
            GRN=8'h61;
            BLU=8'h4F;
        end
        3276:
        begin
            RED=8'h7D;
            GRN=8'h82;
            BLU=8'h6B;
        end
        3277:
        begin
            RED=8'h7C;
            GRN=8'h83;
            BLU=8'h67;
        end
        3278:
        begin
            RED=8'h7C;
            GRN=8'h84;
            BLU=8'h65;
        end
        3279:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h65;
        end
        3280:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h65;
        end
        3281:
        begin
            RED=8'h7F;
            GRN=8'h82;
            BLU=8'h67;
        end
        3282:
        begin
            RED=8'h87;
            GRN=8'h7A;
            BLU=8'h58;
        end
        3283:
        begin
            RED=8'hA9;
            GRN=8'h8E;
            BLU=8'h63;
        end
        3284:
        begin
            RED=8'hCD;
            GRN=8'hAD;
            BLU=8'h78;
        end
        3285:
        begin
            RED=8'hE7;
            GRN=8'hBF;
            BLU=8'h80;
        end
        3286:
        begin
            RED=8'hEE;
            GRN=8'hC1;
            BLU=8'h7E;
        end
        3287:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3288:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3289:
        begin
            RED=8'hEE;
            GRN=8'hC1;
            BLU=8'h80;
        end
        3290:
        begin
            RED=8'hEE;
            GRN=8'hC1;
            BLU=8'h80;
        end
        3291:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3292:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        3293:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        3294:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h82;
        end
        3295:
        begin
            RED=8'hE9;
            GRN=8'hBA;
            BLU=8'h86;
        end
        3296:
        begin
            RED=8'hE1;
            GRN=8'hB3;
            BLU=8'h75;
        end
        3297:
        begin
            RED=8'hEE;
            GRN=8'hC1;
            BLU=8'h80;
        end
        3298:
        begin
            RED=8'hEE;
            GRN=8'hC1;
            BLU=8'h80;
        end
        3299:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3300:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h80;
        end
        3301:
        begin
            RED=8'hEF;
            GRN=8'hBE;
            BLU=8'h82;
        end
        3302:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h82;
        end
        3303:
        begin
            RED=8'hE0;
            GRN=8'hB5;
            BLU=8'h76;
        end
        3304:
        begin
            RED=8'hEA;
            GRN=8'hC0;
            BLU=8'h81;
        end
        3305:
        begin
            RED=8'hF0;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3306:
        begin
            RED=8'hE9;
            GRN=8'hC2;
            BLU=8'h84;
        end
        3307:
        begin
            RED=8'hE0;
            GRN=8'hB8;
            BLU=8'h78;
        end
        3308:
        begin
            RED=8'hE2;
            GRN=8'hBE;
            BLU=8'h88;
        end
        3309:
        begin
            RED=8'hAA;
            GRN=8'h9C;
            BLU=8'h84;
        end
        3310:
        begin
            RED=8'hAD;
            GRN=8'hB3;
            BLU=8'hBA;
        end
        3311:
        begin
            RED=8'hF4;
            GRN=8'hF5;
            BLU=8'hF5;
        end
        3312:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hF9;
        end
        3313:
        begin
            RED=8'hF8;
            GRN=8'hFA;
            BLU=8'hF9;
        end
        3314:
        begin
            RED=8'hE9;
            GRN=8'hEA;
            BLU=8'hE5;
        end
        3315:
        begin
            RED=8'h7A;
            GRN=8'h7C;
            BLU=8'h6C;
        end
        3316:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h68;
        end
        3317:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h63;
        end
        3318:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h64;
        end
        3319:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h65;
        end
        3320:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h63;
        end
        3321:
        begin
            RED=8'h7C;
            GRN=8'h84;
            BLU=8'h67;
        end
        3322:
        begin
            RED=8'h58;
            GRN=8'h61;
            BLU=8'h4C;
        end
        3323:
        begin
            RED=8'h2D;
            GRN=8'h30;
            BLU=8'h25;
        end
        3324:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h28;
        end
        3325:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3326:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3327:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3328:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3329:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3330:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3331:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3332:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3333:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3334:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3335:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h28;
        end
        3336:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3337:
        begin
            RED=8'h30;
            GRN=8'h32;
            BLU=8'h28;
        end
        3338:
        begin
            RED=8'h2C;
            GRN=8'h30;
            BLU=8'h24;
        end
        3339:
        begin
            RED=8'h2C;
            GRN=8'h30;
            BLU=8'h22;
        end
        3340:
        begin
            RED=8'h3F;
            GRN=8'h43;
            BLU=8'h33;
        end
        3341:
        begin
            RED=8'h70;
            GRN=8'h75;
            BLU=8'h61;
        end
        3342:
        begin
            RED=8'h7C;
            GRN=8'h85;
            BLU=8'h65;
        end
        3343:
        begin
            RED=8'h7D;
            GRN=8'h83;
            BLU=8'h66;
        end
        3344:
        begin
            RED=8'h7F;
            GRN=8'h82;
            BLU=8'h69;
        end
        3345:
        begin
            RED=8'h82;
            GRN=8'h84;
            BLU=8'h6D;
        end
        3346:
        begin
            RED=8'h7F;
            GRN=8'h82;
            BLU=8'h6B;
        end
        3347:
        begin
            RED=8'h82;
            GRN=8'h83;
            BLU=8'h68;
        end
        3348:
        begin
            RED=8'h80;
            GRN=8'h77;
            BLU=8'h51;
        end
        3349:
        begin
            RED=8'hD8;
            GRN=8'hBB;
            BLU=8'h86;
        end
        3350:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        3351:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3352:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3353:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3354:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3355:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        3356:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        3357:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        3358:
        begin
            RED=8'hEC;
            GRN=8'hBE;
            BLU=8'h7F;
        end
        3359:
        begin
            RED=8'hEF;
            GRN=8'hC1;
            BLU=8'h84;
        end
        3360:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h7F;
        end
        3361:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3362:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3363:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3364:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h80;
        end
        3365:
        begin
            RED=8'hEF;
            GRN=8'hBE;
            BLU=8'h83;
        end
        3366:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h84;
        end
        3367:
        begin
            RED=8'hDE;
            GRN=8'hB1;
            BLU=8'h77;
        end
        3368:
        begin
            RED=8'hDF;
            GRN=8'hB3;
            BLU=8'h7C;
        end
        3369:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h81;
        end
        3370:
        begin
            RED=8'hE8;
            GRN=8'hC2;
            BLU=8'h82;
        end
        3371:
        begin
            RED=8'hDB;
            GRN=8'hB3;
            BLU=8'h72;
        end
        3372:
        begin
            RED=8'hD0;
            GRN=8'hB0;
            BLU=8'h85;
        end
        3373:
        begin
            RED=8'hA5;
            GRN=8'hA0;
            BLU=8'h98;
        end
        3374:
        begin
            RED=8'hCA;
            GRN=8'hD5;
            BLU=8'hE2;
        end
        3375:
        begin
            RED=8'hC7;
            GRN=8'hCA;
            BLU=8'hD0;
        end
        3376:
        begin
            RED=8'hFC;
            GRN=8'hFB;
            BLU=8'hFC;
        end
        3377:
        begin
            RED=8'hFA;
            GRN=8'hFB;
            BLU=8'hFB;
        end
        3378:
        begin
            RED=8'hF8;
            GRN=8'hF9;
            BLU=8'hF9;
        end
        3379:
        begin
            RED=8'hCD;
            GRN=8'hCE;
            BLU=8'hC9;
        end
        3380:
        begin
            RED=8'h77;
            GRN=8'h7A;
            BLU=8'h6A;
        end
        3381:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h69;
        end
        3382:
        begin
            RED=8'h7F;
            GRN=8'h84;
            BLU=8'h63;
        end
        3383:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h65;
        end
        3384:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h63;
        end
        3385:
        begin
            RED=8'h7B;
            GRN=8'h84;
            BLU=8'h66;
        end
        3386:
        begin
            RED=8'h58;
            GRN=8'h61;
            BLU=8'h4C;
        end
        3387:
        begin
            RED=8'h2D;
            GRN=8'h31;
            BLU=8'h25;
        end
        3388:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h28;
        end
        3389:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3390:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3391:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3392:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3393:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3394:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3395:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3396:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3397:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3398:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3399:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3400:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3401:
        begin
            RED=8'h2F;
            GRN=8'h32;
            BLU=8'h29;
        end
        3402:
        begin
            RED=8'h2F;
            GRN=8'h32;
            BLU=8'h29;
        end
        3403:
        begin
            RED=8'h2E;
            GRN=8'h31;
            BLU=8'h28;
        end
        3404:
        begin
            RED=8'h2C;
            GRN=8'h2F;
            BLU=8'h26;
        end
        3405:
        begin
            RED=8'h2D;
            GRN=8'h31;
            BLU=8'h26;
        end
        3406:
        begin
            RED=8'h5A;
            GRN=8'h60;
            BLU=8'h4C;
        end
        3407:
        begin
            RED=8'h7C;
            GRN=8'h80;
            BLU=8'h6A;
        end
        3408:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h69;
        end
        3409:
        begin
            RED=8'h7F;
            GRN=8'h82;
            BLU=8'h66;
        end
        3410:
        begin
            RED=8'h7D;
            GRN=8'h83;
            BLU=8'h66;
        end
        3411:
        begin
            RED=8'h7A;
            GRN=8'h84;
            BLU=8'h69;
        end
        3412:
        begin
            RED=8'h7E;
            GRN=8'h82;
            BLU=8'h64;
        end
        3413:
        begin
            RED=8'h8B;
            GRN=8'h7E;
            BLU=8'h54;
        end
        3414:
        begin
            RED=8'hE0;
            GRN=8'hBE;
            BLU=8'h88;
        end
        3415:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        3416:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3417:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3418:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3419:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        3420:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7C;
        end
        3421:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h80;
        end
        3422:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3423:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7B;
        end
        3424:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        3425:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3426:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3427:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3428:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        3429:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        3430:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h80;
        end
        3431:
        begin
            RED=8'hEC;
            GRN=8'hBF;
            BLU=8'h85;
        end
        3432:
        begin
            RED=8'hC6;
            GRN=8'h9C;
            BLU=8'h64;
        end
        3433:
        begin
            RED=8'hE7;
            GRN=8'hBD;
            BLU=8'h81;
        end
        3434:
        begin
            RED=8'hE8;
            GRN=8'hC3;
            BLU=8'h81;
        end
        3435:
        begin
            RED=8'hEA;
            GRN=8'hC3;
            BLU=8'h7F;
        end
        3436:
        begin
            RED=8'hB3;
            GRN=8'h97;
            BLU=8'h76;
        end
        3437:
        begin
            RED=8'hB6;
            GRN=8'hB7;
            BLU=8'hC4;
        end
        3438:
        begin
            RED=8'hD2;
            GRN=8'hE0;
            BLU=8'hF4;
        end
        3439:
        begin
            RED=8'hA3;
            GRN=8'hA8;
            BLU=8'hB3;
        end
        3440:
        begin
            RED=8'hFA;
            GRN=8'hFA;
            BLU=8'hFD;
        end
        3441:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFE;
        end
        3442:
        begin
            RED=8'hFA;
            GRN=8'hFA;
            BLU=8'hFA;
        end
        3443:
        begin
            RED=8'hF7;
            GRN=8'hF7;
            BLU=8'hF7;
        end
        3444:
        begin
            RED=8'h85;
            GRN=8'h86;
            BLU=8'h81;
        end
        3445:
        begin
            RED=8'h77;
            GRN=8'h7A;
            BLU=8'h6A;
        end
        3446:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h68;
        end
        3447:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h65;
        end
        3448:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h63;
        end
        3449:
        begin
            RED=8'h7B;
            GRN=8'h84;
            BLU=8'h66;
        end
        3450:
        begin
            RED=8'h58;
            GRN=8'h61;
            BLU=8'h4C;
        end
        3451:
        begin
            RED=8'h2D;
            GRN=8'h30;
            BLU=8'h25;
        end
        3452:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h28;
        end
        3453:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3454:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3455:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3456:
        begin
            RED=8'h2F;
            GRN=8'h2F;
            BLU=8'h25;
        end
        3457:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h28;
        end
        3458:
        begin
            RED=8'h31;
            GRN=8'h31;
            BLU=8'h2A;
        end
        3459:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3460:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3461:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3462:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3463:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3464:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3465:
        begin
            RED=8'h2F;
            GRN=8'h32;
            BLU=8'h29;
        end
        3466:
        begin
            RED=8'h2F;
            GRN=8'h32;
            BLU=8'h29;
        end
        3467:
        begin
            RED=8'h30;
            GRN=8'h33;
            BLU=8'h2C;
        end
        3468:
        begin
            RED=8'h2E;
            GRN=8'h30;
            BLU=8'h2A;
        end
        3469:
        begin
            RED=8'h2F;
            GRN=8'h31;
            BLU=8'h2C;
        end
        3470:
        begin
            RED=8'h2C;
            GRN=8'h2F;
            BLU=8'h26;
        end
        3471:
        begin
            RED=8'h3F;
            GRN=8'h43;
            BLU=8'h33;
        end
        3472:
        begin
            RED=8'h76;
            GRN=8'h79;
            BLU=8'h61;
        end
        3473:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h62;
        end
        3474:
        begin
            RED=8'h81;
            GRN=8'h83;
            BLU=8'h5D;
        end
        3475:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h60;
        end
        3476:
        begin
            RED=8'h7C;
            GRN=8'h84;
            BLU=8'h67;
        end
        3477:
        begin
            RED=8'h81;
            GRN=8'h80;
            BLU=8'h5F;
        end
        3478:
        begin
            RED=8'h91;
            GRN=8'h7F;
            BLU=8'h54;
        end
        3479:
        begin
            RED=8'hDF;
            GRN=8'hB8;
            BLU=8'h7D;
        end
        3480:
        begin
            RED=8'hEA;
            GRN=8'hC0;
            BLU=8'h81;
        end
        3481:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3482:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        3483:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7B;
        end
        3484:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        3485:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h82;
        end
        3486:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3487:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h78;
        end
        3488:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        3489:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h80;
        end
        3490:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3491:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3492:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        3493:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h79;
        end
        3494:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h7B;
        end
        3495:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h80;
        end
        3496:
        begin
            RED=8'hE8;
            GRN=8'hBD;
            BLU=8'h84;
        end
        3497:
        begin
            RED=8'hC6;
            GRN=8'h9D;
            BLU=8'h63;
        end
        3498:
        begin
            RED=8'hE6;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3499:
        begin
            RED=8'hEB;
            GRN=8'hC4;
            BLU=8'h82;
        end
        3500:
        begin
            RED=8'hAD;
            GRN=8'h98;
            BLU=8'h80;
        end
        3501:
        begin
            RED=8'hCF;
            GRN=8'hD7;
            BLU=8'hEF;
        end
        3502:
        begin
            RED=8'hD0;
            GRN=8'hE0;
            BLU=8'hF9;
        end
        3503:
        begin
            RED=8'hB7;
            GRN=8'hBE;
            BLU=8'hCD;
        end
        3504:
        begin
            RED=8'hF1;
            GRN=8'hF2;
            BLU=8'hF6;
        end
        3505:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFE;
        end
        3506:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hF9;
        end
        3507:
        begin
            RED=8'hFA;
            GRN=8'hFA;
            BLU=8'hF9;
        end
        3508:
        begin
            RED=8'hE0;
            GRN=8'hE0;
            BLU=8'hE1;
        end
        3509:
        begin
            RED=8'hAD;
            GRN=8'hAE;
            BLU=8'hA8;
        end
        3510:
        begin
            RED=8'h77;
            GRN=8'h7A;
            BLU=8'h6B;
        end
        3511:
        begin
            RED=8'h7D;
            GRN=8'h81;
            BLU=8'h67;
        end
        3512:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h64;
        end
        3513:
        begin
            RED=8'h7C;
            GRN=8'h84;
            BLU=8'h66;
        end
        3514:
        begin
            RED=8'h58;
            GRN=8'h61;
            BLU=8'h4C;
        end
        3515:
        begin
            RED=8'h2D;
            GRN=8'h30;
            BLU=8'h25;
        end
        3516:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h28;
        end
        3517:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3518:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3519:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3520:
        begin
            RED=8'h68;
            GRN=8'h66;
            BLU=8'h53;
        end
        3521:
        begin
            RED=8'h36;
            GRN=8'h33;
            BLU=8'h27;
        end
        3522:
        begin
            RED=8'h31;
            GRN=8'h2F;
            BLU=8'h2B;
        end
        3523:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h2C;
        end
        3524:
        begin
            RED=8'h32;
            GRN=8'h33;
            BLU=8'h2B;
        end
        3525:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3526:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3527:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3528:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3529:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3530:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3531:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3532:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3533:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3534:
        begin
            RED=8'h2E;
            GRN=8'h2F;
            BLU=8'h29;
        end
        3535:
        begin
            RED=8'h2E;
            GRN=8'h30;
            BLU=8'h25;
        end
        3536:
        begin
            RED=8'h30;
            GRN=8'h32;
            BLU=8'h23;
        end
        3537:
        begin
            RED=8'h60;
            GRN=8'h63;
            BLU=8'h4E;
        end
        3538:
        begin
            RED=8'h7C;
            GRN=8'h81;
            BLU=8'h64;
        end
        3539:
        begin
            RED=8'h7E;
            GRN=8'h84;
            BLU=8'h64;
        end
        3540:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h62;
        end
        3541:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h61;
        end
        3542:
        begin
            RED=8'h7E;
            GRN=8'h83;
            BLU=8'h5F;
        end
        3543:
        begin
            RED=8'h87;
            GRN=8'h7D;
            BLU=8'h55;
        end
        3544:
        begin
            RED=8'hB4;
            GRN=8'hA2;
            BLU=8'h6F;
        end
        3545:
        begin
            RED=8'hDF;
            GRN=8'hC2;
            BLU=8'h84;
        end
        3546:
        begin
            RED=8'hED;
            GRN=8'hC3;
            BLU=8'h82;
        end
        3547:
        begin
            RED=8'hED;
            GRN=8'hBF;
            BLU=8'h7F;
        end
        3548:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h81;
        end
        3549:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h80;
        end
        3550:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h7F;
        end
        3551:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3552:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h81;
        end
        3553:
        begin
            RED=8'hEE;
            GRN=8'hC2;
            BLU=8'h81;
        end
        3554:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7E;
        end
        3555:
        begin
            RED=8'hEE;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        3556:
        begin
            RED=8'hEE;
            GRN=8'hBF;
            BLU=8'h7E;
        end
        3557:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h80;
        end
        3558:
        begin
            RED=8'hEC;
            GRN=8'hC1;
            BLU=8'h7D;
        end
        3559:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h7C;
        end
        3560:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        3561:
        begin
            RED=8'hE6;
            GRN=8'hB8;
            BLU=8'h81;
        end
        3562:
        begin
            RED=8'hD3;
            GRN=8'hA6;
            BLU=8'h72;
        end
        3563:
        begin
            RED=8'hD7;
            GRN=8'hB7;
            BLU=8'h90;
        end
        3564:
        begin
            RED=8'hBE;
            GRN=8'hBD;
            BLU=8'hB9;
        end
        3565:
        begin
            RED=8'hCC;
            GRN=8'hE0;
            BLU=8'hFA;
        end
        3566:
        begin
            RED=8'hD1;
            GRN=8'hE0;
            BLU=8'hFC;
        end
        3567:
        begin
            RED=8'hC6;
            GRN=8'hD2;
            BLU=8'hE0;
        end
        3568:
        begin
            RED=8'hE2;
            GRN=8'hE8;
            BLU=8'hEB;
        end
        3569:
        begin
            RED=8'hFB;
            GRN=8'hFD;
            BLU=8'hFC;
        end
        3570:
        begin
            RED=8'hFD;
            GRN=8'hFD;
            BLU=8'hFC;
        end
        3571:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        3572:
        begin
            RED=8'hF7;
            GRN=8'hF7;
            BLU=8'hF7;
        end
        3573:
        begin
            RED=8'hC4;
            GRN=8'hC4;
            BLU=8'hC4;
        end
        3574:
        begin
            RED=8'hE9;
            GRN=8'hEA;
            BLU=8'hE9;
        end
        3575:
        begin
            RED=8'h93;
            GRN=8'h96;
            BLU=8'h8D;
        end
        3576:
        begin
            RED=8'h78;
            GRN=8'h7E;
            BLU=8'h67;
        end
        3577:
        begin
            RED=8'h7F;
            GRN=8'h85;
            BLU=8'h68;
        end
        3578:
        begin
            RED=8'h5F;
            GRN=8'h63;
            BLU=8'h51;
        end
        3579:
        begin
            RED=8'h2E;
            GRN=8'h2F;
            BLU=8'h26;
        end
        3580:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h28;
        end
        3581:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3582:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3583:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3584:
        begin
            RED=8'hB5;
            GRN=8'hB3;
            BLU=8'h9E;
        end
        3585:
        begin
            RED=8'h4F;
            GRN=8'h4D;
            BLU=8'h40;
        end
        3586:
        begin
            RED=8'h27;
            GRN=8'h25;
            BLU=8'h20;
        end
        3587:
        begin
            RED=8'h2D;
            GRN=8'h2E;
            BLU=8'h29;
        end
        3588:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3589:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3590:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3591:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3592:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3593:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3594:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3595:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3596:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3597:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3598:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h2B;
        end
        3599:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h28;
        end
        3600:
        begin
            RED=8'h31;
            GRN=8'h33;
            BLU=8'h25;
        end
        3601:
        begin
            RED=8'h2E;
            GRN=8'h31;
            BLU=8'h20;
        end
        3602:
        begin
            RED=8'h47;
            GRN=8'h4B;
            BLU=8'h36;
        end
        3603:
        begin
            RED=8'h76;
            GRN=8'h7C;
            BLU=8'h62;
        end
        3604:
        begin
            RED=8'h7E;
            GRN=8'h84;
            BLU=8'h66;
        end
        3605:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h64;
        end
        3606:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h63;
        end
        3607:
        begin
            RED=8'h7F;
            GRN=8'h84;
            BLU=8'h61;
        end
        3608:
        begin
            RED=8'h83;
            GRN=8'h82;
            BLU=8'h58;
        end
        3609:
        begin
            RED=8'h89;
            GRN=8'h80;
            BLU=8'h4F;
        end
        3610:
        begin
            RED=8'hB3;
            GRN=8'hA0;
            BLU=8'h70;
        end
        3611:
        begin
            RED=8'hDC;
            GRN=8'hBD;
            BLU=8'h90;
        end
        3612:
        begin
            RED=8'hE9;
            GRN=8'hC0;
            BLU=8'h8A;
        end
        3613:
        begin
            RED=8'hEA;
            GRN=8'hC2;
            BLU=8'h7D;
        end
        3614:
        begin
            RED=8'hED;
            GRN=8'hC1;
            BLU=8'h7A;
        end
        3615:
        begin
            RED=8'hEF;
            GRN=8'hBF;
            BLU=8'h7F;
        end
        3616:
        begin
            RED=8'hEA;
            GRN=8'hBD;
            BLU=8'h7D;
        end
        3617:
        begin
            RED=8'hE6;
            GRN=8'hBA;
            BLU=8'h79;
        end
        3618:
        begin
            RED=8'hE1;
            GRN=8'hB5;
            BLU=8'h75;
        end
        3619:
        begin
            RED=8'hEB;
            GRN=8'hC0;
            BLU=8'h80;
        end
        3620:
        begin
            RED=8'hEC;
            GRN=8'hC1;
            BLU=8'h80;
        end
        3621:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3622:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h81;
        end
        3623:
        begin
            RED=8'hE9;
            GRN=8'hC2;
            BLU=8'h7F;
        end
        3624:
        begin
            RED=8'hE7;
            GRN=8'hC3;
            BLU=8'h7B;
        end
        3625:
        begin
            RED=8'hE7;
            GRN=8'hBD;
            BLU=8'h8B;
        end
        3626:
        begin
            RED=8'hBC;
            GRN=8'hA1;
            BLU=8'h81;
        end
        3627:
        begin
            RED=8'hAF;
            GRN=8'hA9;
            BLU=8'hA2;
        end
        3628:
        begin
            RED=8'hD2;
            GRN=8'hDA;
            BLU=8'hED;
        end
        3629:
        begin
            RED=8'hD0;
            GRN=8'hDF;
            BLU=8'hFE;
        end
        3630:
        begin
            RED=8'hD1;
            GRN=8'hDE;
            BLU=8'hFB;
        end
        3631:
        begin
            RED=8'hCE;
            GRN=8'hD9;
            BLU=8'hE7;
        end
        3632:
        begin
            RED=8'hD3;
            GRN=8'hD9;
            BLU=8'hDC;
        end
        3633:
        begin
            RED=8'hFA;
            GRN=8'hFC;
            BLU=8'hFB;
        end
        3634:
        begin
            RED=8'hFD;
            GRN=8'hFD;
            BLU=8'hFC;
        end
        3635:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        3636:
        begin
            RED=8'hFA;
            GRN=8'hFA;
            BLU=8'hFA;
        end
        3637:
        begin
            RED=8'hC9;
            GRN=8'hC9;
            BLU=8'hC9;
        end
        3638:
        begin
            RED=8'hF7;
            GRN=8'hF7;
            BLU=8'hF7;
        end
        3639:
        begin
            RED=8'hF6;
            GRN=8'hF8;
            BLU=8'hF3;
        end
        3640:
        begin
            RED=8'hB7;
            GRN=8'hBB;
            BLU=8'hAB;
        end
        3641:
        begin
            RED=8'h71;
            GRN=8'h75;
            BLU=8'h61;
        end
        3642:
        begin
            RED=8'h5D;
            GRN=8'h60;
            BLU=8'h53;
        end
        3643:
        begin
            RED=8'h2E;
            GRN=8'h30;
            BLU=8'h28;
        end
        3644:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h28;
        end
        3645:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3646:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3647:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3648:
        begin
            RED=8'hB2;
            GRN=8'hB0;
            BLU=8'h9C;
        end
        3649:
        begin
            RED=8'h50;
            GRN=8'h4D;
            BLU=8'h41;
        end
        3650:
        begin
            RED=8'h31;
            GRN=8'h2F;
            BLU=8'h2A;
        end
        3651:
        begin
            RED=8'h2A;
            GRN=8'h2B;
            BLU=8'h25;
        end
        3652:
        begin
            RED=8'h27;
            GRN=8'h28;
            BLU=8'h20;
        end
        3653:
        begin
            RED=8'h2E;
            GRN=8'h2F;
            BLU=8'h27;
        end
        3654:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3655:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h28;
        end
        3656:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3657:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3658:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3659:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3660:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3661:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3662:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3663:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3664:
        begin
            RED=8'h30;
            GRN=8'h32;
            BLU=8'h27;
        end
        3665:
        begin
            RED=8'h30;
            GRN=8'h32;
            BLU=8'h26;
        end
        3666:
        begin
            RED=8'h2E;
            GRN=8'h31;
            BLU=8'h24;
        end
        3667:
        begin
            RED=8'h33;
            GRN=8'h37;
            BLU=8'h28;
        end
        3668:
        begin
            RED=8'h6E;
            GRN=8'h73;
            BLU=8'h5F;
        end
        3669:
        begin
            RED=8'h7C;
            GRN=8'h82;
            BLU=8'h67;
        end
        3670:
        begin
            RED=8'h7E;
            GRN=8'h86;
            BLU=8'h68;
        end
        3671:
        begin
            RED=8'h79;
            GRN=8'h85;
            BLU=8'h67;
        end
        3672:
        begin
            RED=8'h7B;
            GRN=8'h85;
            BLU=8'h63;
        end
        3673:
        begin
            RED=8'h7F;
            GRN=8'h83;
            BLU=8'h63;
        end
        3674:
        begin
            RED=8'h7B;
            GRN=8'h7A;
            BLU=8'h61;
        end
        3675:
        begin
            RED=8'hBE;
            GRN=8'hB3;
            BLU=8'h97;
        end
        3676:
        begin
            RED=8'hC2;
            GRN=8'hAB;
            BLU=8'h80;
        end
        3677:
        begin
            RED=8'hDB;
            GRN=8'hBE;
            BLU=8'h85;
        end
        3678:
        begin
            RED=8'hE6;
            GRN=8'hC2;
            BLU=8'h80;
        end
        3679:
        begin
            RED=8'hEB;
            GRN=8'hC1;
            BLU=8'h7A;
        end
        3680:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        3681:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3682:
        begin
            RED=8'hD1;
            GRN=8'hA8;
            BLU=8'h69;
        end
        3683:
        begin
            RED=8'hD3;
            GRN=8'hAD;
            BLU=8'h70;
        end
        3684:
        begin
            RED=8'hEB;
            GRN=8'hC4;
            BLU=8'h88;
        end
        3685:
        begin
            RED=8'hEC;
            GRN=8'hC2;
            BLU=8'h80;
        end
        3686:
        begin
            RED=8'hE7;
            GRN=8'hC4;
            BLU=8'h84;
        end
        3687:
        begin
            RED=8'hCA;
            GRN=8'hAA;
            BLU=8'h8C;
        end
        3688:
        begin
            RED=8'h74;
            GRN=8'h55;
            BLU=8'h64;
        end
        3689:
        begin
            RED=8'h4E;
            GRN=8'h25;
            BLU=8'h4F;
        end
        3690:
        begin
            RED=8'h41;
            GRN=8'h2B;
            BLU=8'h58;
        end
        3691:
        begin
            RED=8'hAA;
            GRN=8'hB0;
            BLU=8'hD5;
        end
        3692:
        begin
            RED=8'hCE;
            GRN=8'hDE;
            BLU=8'hFB;
        end
        3693:
        begin
            RED=8'hD2;
            GRN=8'hDF;
            BLU=8'hF9;
        end
        3694:
        begin
            RED=8'hD0;
            GRN=8'hDD;
            BLU=8'hFA;
        end
        3695:
        begin
            RED=8'hCC;
            GRN=8'hD7;
            BLU=8'hE5;
        end
        3696:
        begin
            RED=8'hCF;
            GRN=8'hD4;
            BLU=8'hD7;
        end
        3697:
        begin
            RED=8'hFC;
            GRN=8'hFD;
            BLU=8'hFD;
        end
        3698:
        begin
            RED=8'hFB;
            GRN=8'hFB;
            BLU=8'hFB;
        end
        3699:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        3700:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        3701:
        begin
            RED=8'hD8;
            GRN=8'hD8;
            BLU=8'hD8;
        end
        3702:
        begin
            RED=8'hF2;
            GRN=8'hF2;
            BLU=8'hF2;
        end
        3703:
        begin
            RED=8'hFB;
            GRN=8'hFD;
            BLU=8'hFC;
        end
        3704:
        begin
            RED=8'hFA;
            GRN=8'hFC;
            BLU=8'hF6;
        end
        3705:
        begin
            RED=8'hD8;
            GRN=8'hDA;
            BLU=8'hD1;
        end
        3706:
        begin
            RED=8'h5B;
            GRN=8'h5E;
            BLU=8'h57;
        end
        3707:
        begin
            RED=8'h2E;
            GRN=8'h30;
            BLU=8'h28;
        end
        3708:
        begin
            RED=8'h2E;
            GRN=8'h2F;
            BLU=8'h27;
        end
        3709:
        begin
            RED=8'h31;
            GRN=8'h32;
            BLU=8'h2A;
        end
        3710:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3711:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3712:
        begin
            RED=8'hB2;
            GRN=8'hB0;
            BLU=8'h9C;
        end
        3713:
        begin
            RED=8'h50;
            GRN=8'h4D;
            BLU=8'h41;
        end
        3714:
        begin
            RED=8'h33;
            GRN=8'h31;
            BLU=8'h2C;
        end
        3715:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h2C;
        end
        3716:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h2A;
        end
        3717:
        begin
            RED=8'h2A;
            GRN=8'h2B;
            BLU=8'h23;
        end
        3718:
        begin
            RED=8'h2A;
            GRN=8'h2B;
            BLU=8'h23;
        end
        3719:
        begin
            RED=8'h2D;
            GRN=8'h2E;
            BLU=8'h26;
        end
        3720:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h28;
        end
        3721:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3722:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3723:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3724:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3725:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3726:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3727:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3728:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h2B;
        end
        3729:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h2B;
        end
        3730:
        begin
            RED=8'h2F;
            GRN=8'h31;
            BLU=8'h2C;
        end
        3731:
        begin
            RED=8'h2D;
            GRN=8'h30;
            BLU=8'h2A;
        end
        3732:
        begin
            RED=8'h2D;
            GRN=8'h31;
            BLU=8'h24;
        end
        3733:
        begin
            RED=8'h61;
            GRN=8'h65;
            BLU=8'h50;
        end
        3734:
        begin
            RED=8'h7C;
            GRN=8'h83;
            BLU=8'h67;
        end
        3735:
        begin
            RED=8'h7D;
            GRN=8'h84;
            BLU=8'h6A;
        end
        3736:
        begin
            RED=8'h7E;
            GRN=8'h85;
            BLU=8'h6A;
        end
        3737:
        begin
            RED=8'h7D;
            GRN=8'h82;
            BLU=8'h6D;
        end
        3738:
        begin
            RED=8'hB1;
            GRN=8'hB3;
            BLU=8'hAB;
        end
        3739:
        begin
            RED=8'hF7;
            GRN=8'hF7;
            BLU=8'hF0;
        end
        3740:
        begin
            RED=8'hF0;
            GRN=8'hE9;
            BLU=8'hE5;
        end
        3741:
        begin
            RED=8'hB2;
            GRN=8'hA0;
            BLU=8'hA2;
        end
        3742:
        begin
            RED=8'hAE;
            GRN=8'h90;
            BLU=8'h7D;
        end
        3743:
        begin
            RED=8'hE2;
            GRN=8'hC1;
            BLU=8'h88;
        end
        3744:
        begin
            RED=8'hED;
            GRN=8'hC0;
            BLU=8'h7D;
        end
        3745:
        begin
            RED=8'hEC;
            GRN=8'hC0;
            BLU=8'h7F;
        end
        3746:
        begin
            RED=8'hE9;
            GRN=8'hC1;
            BLU=8'h85;
        end
        3747:
        begin
            RED=8'hDA;
            GRN=8'hB7;
            BLU=8'h7D;
        end
        3748:
        begin
            RED=8'hC6;
            GRN=8'hA5;
            BLU=8'h6B;
        end
        3749:
        begin
            RED=8'hE2;
            GRN=8'hBD;
            BLU=8'h91;
        end
        3750:
        begin
            RED=8'h95;
            GRN=8'h73;
            BLU=8'h76;
        end
        3751:
        begin
            RED=8'h3E;
            GRN=8'h21;
            BLU=8'h57;
        end
        3752:
        begin
            RED=8'h37;
            GRN=8'h1F;
            BLU=8'h75;
        end
        3753:
        begin
            RED=8'h3A;
            GRN=8'h1B;
            BLU=8'h7E;
        end
        3754:
        begin
            RED=8'h38;
            GRN=8'h22;
            BLU=8'h76;
        end
        3755:
        begin
            RED=8'h45;
            GRN=8'h43;
            BLU=8'h79;
        end
        3756:
        begin
            RED=8'hCD;
            GRN=8'hDB;
            BLU=8'hF8;
        end
        3757:
        begin
            RED=8'hCF;
            GRN=8'hE2;
            BLU=8'hF9;
        end
        3758:
        begin
            RED=8'hD1;
            GRN=8'hDF;
            BLU=8'hFC;
        end
        3759:
        begin
            RED=8'hCA;
            GRN=8'hD5;
            BLU=8'hE3;
        end
        3760:
        begin
            RED=8'hDE;
            GRN=8'hE4;
            BLU=8'hE7;
        end
        3761:
        begin
            RED=8'hFC;
            GRN=8'hFE;
            BLU=8'hFD;
        end
        3762:
        begin
            RED=8'hFB;
            GRN=8'hFB;
            BLU=8'hFB;
        end
        3763:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        3764:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        3765:
        begin
            RED=8'hDC;
            GRN=8'hDC;
            BLU=8'hDC;
        end
        3766:
        begin
            RED=8'hF4;
            GRN=8'hF4;
            BLU=8'hF4;
        end
        3767:
        begin
            RED=8'hFC;
            GRN=8'hFD;
            BLU=8'hFF;
        end
        3768:
        begin
            RED=8'hFA;
            GRN=8'hFB;
            BLU=8'hFE;
        end
        3769:
        begin
            RED=8'hF9;
            GRN=8'hFB;
            BLU=8'hFB;
        end
        3770:
        begin
            RED=8'hE2;
            GRN=8'hE4;
            BLU=8'hE1;
        end
        3771:
        begin
            RED=8'h54;
            GRN=8'h56;
            BLU=8'h4F;
        end
        3772:
        begin
            RED=8'h2D;
            GRN=8'h2E;
            BLU=8'h26;
        end
        3773:
        begin
            RED=8'h2E;
            GRN=8'h2F;
            BLU=8'h27;
        end
        3774:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3775:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3776:
        begin
            RED=8'hB2;
            GRN=8'hB0;
            BLU=8'hA0;
        end
        3777:
        begin
            RED=8'h51;
            GRN=8'h50;
            BLU=8'h43;
        end
        3778:
        begin
            RED=8'h32;
            GRN=8'h31;
            BLU=8'h26;
        end
        3779:
        begin
            RED=8'h32;
            GRN=8'h32;
            BLU=8'h28;
        end
        3780:
        begin
            RED=8'h31;
            GRN=8'h32;
            BLU=8'h27;
        end
        3781:
        begin
            RED=8'h31;
            GRN=8'h32;
            BLU=8'h28;
        end
        3782:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h27;
        end
        3783:
        begin
            RED=8'h28;
            GRN=8'h29;
            BLU=8'h21;
        end
        3784:
        begin
            RED=8'h2E;
            GRN=8'h2F;
            BLU=8'h29;
        end
        3785:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3786:
        begin
            RED=8'h31;
            GRN=8'h32;
            BLU=8'h2A;
        end
        3787:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3788:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3789:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3790:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3791:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3792:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h2A;
        end
        3793:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h2A;
        end
        3794:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h2B;
        end
        3795:
        begin
            RED=8'h2F;
            GRN=8'h31;
            BLU=8'h2A;
        end
        3796:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h27;
        end
        3797:
        begin
            RED=8'h30;
            GRN=8'h32;
            BLU=8'h25;
        end
        3798:
        begin
            RED=8'h47;
            GRN=8'h4A;
            BLU=8'h3A;
        end
        3799:
        begin
            RED=8'h7C;
            GRN=8'h7F;
            BLU=8'h68;
        end
        3800:
        begin
            RED=8'h7F;
            GRN=8'h82;
            BLU=8'h6E;
        end
        3801:
        begin
            RED=8'h7B;
            GRN=8'h7D;
            BLU=8'h6F;
        end
        3802:
        begin
            RED=8'hF2;
            GRN=8'hF2;
            BLU=8'hEE;
        end
        3803:
        begin
            RED=8'hF1;
            GRN=8'hF0;
            BLU=8'hF2;
        end
        3804:
        begin
            RED=8'h62;
            GRN=8'h56;
            BLU=8'h81;
        end
        3805:
        begin
            RED=8'h36;
            GRN=8'h20;
            BLU=8'h67;
        end
        3806:
        begin
            RED=8'h38;
            GRN=8'h1E;
            BLU=8'h53;
        end
        3807:
        begin
            RED=8'h6D;
            GRN=8'h53;
            BLU=8'h5D;
        end
        3808:
        begin
            RED=8'hE2;
            GRN=8'hBC;
            BLU=8'h88;
        end
        3809:
        begin
            RED=8'hEA;
            GRN=8'hC3;
            BLU=8'h86;
        end
        3810:
        begin
            RED=8'hE7;
            GRN=8'hC3;
            BLU=8'h85;
        end
        3811:
        begin
            RED=8'hE3;
            GRN=8'hC1;
            BLU=8'h85;
        end
        3812:
        begin
            RED=8'hCD;
            GRN=8'hB0;
            BLU=8'h84;
        end
        3813:
        begin
            RED=8'h74;
            GRN=8'h5C;
            BLU=8'h66;
        end
        3814:
        begin
            RED=8'h3D;
            GRN=8'h20;
            BLU=8'h66;
        end
        3815:
        begin
            RED=8'h38;
            GRN=8'h1D;
            BLU=8'h7F;
        end
        3816:
        begin
            RED=8'h36;
            GRN=8'h20;
            BLU=8'h78;
        end
        3817:
        begin
            RED=8'h37;
            GRN=8'h1D;
            BLU=8'h7A;
        end
        3818:
        begin
            RED=8'h35;
            GRN=8'h1E;
            BLU=8'h75;
        end
        3819:
        begin
            RED=8'h3B;
            GRN=8'h34;
            BLU=8'h6B;
        end
        3820:
        begin
            RED=8'hCD;
            GRN=8'hD6;
            BLU=8'hF4;
        end
        3821:
        begin
            RED=8'hCF;
            GRN=8'hE0;
            BLU=8'hFD;
        end
        3822:
        begin
            RED=8'hD2;
            GRN=8'hE0;
            BLU=8'hFC;
        end
        3823:
        begin
            RED=8'hC3;
            GRN=8'hCB;
            BLU=8'hDA;
        end
        3824:
        begin
            RED=8'hEC;
            GRN=8'hED;
            BLU=8'hF2;
        end
        3825:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFE;
        end
        3826:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        3827:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        3828:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        3829:
        begin
            RED=8'hDD;
            GRN=8'hDD;
            BLU=8'hDD;
        end
        3830:
        begin
            RED=8'hF3;
            GRN=8'hF3;
            BLU=8'hF3;
        end
        3831:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFD;
        end
        3832:
        begin
            RED=8'hFB;
            GRN=8'hFC;
            BLU=8'hFE;
        end
        3833:
        begin
            RED=8'hFB;
            GRN=8'hFB;
            BLU=8'hFC;
        end
        3834:
        begin
            RED=8'hFA;
            GRN=8'hFA;
            BLU=8'hFA;
        end
        3835:
        begin
            RED=8'hEB;
            GRN=8'hEC;
            BLU=8'hE9;
        end
        3836:
        begin
            RED=8'h4F;
            GRN=8'h50;
            BLU=8'h4B;
        end
        3837:
        begin
            RED=8'h2E;
            GRN=8'h2F;
            BLU=8'h28;
        end
        3838:
        begin
            RED=8'h2E;
            GRN=8'h2F;
            BLU=8'h27;
        end
        3839:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3840:
        begin
            RED=8'hAC;
            GRN=8'hA8;
            BLU=8'h96;
        end
        3841:
        begin
            RED=8'h7D;
            GRN=8'h79;
            BLU=8'h66;
        end
        3842:
        begin
            RED=8'h6E;
            GRN=8'h6A;
            BLU=8'h58;
        end
        3843:
        begin
            RED=8'h6E;
            GRN=8'h6A;
            BLU=8'h57;
        end
        3844:
        begin
            RED=8'h6E;
            GRN=8'h69;
            BLU=8'h57;
        end
        3845:
        begin
            RED=8'h6B;
            GRN=8'h69;
            BLU=8'h58;
        end
        3846:
        begin
            RED=8'h6B;
            GRN=8'h69;
            BLU=8'h5A;
        end
        3847:
        begin
            RED=8'h68;
            GRN=8'h66;
            BLU=8'h59;
        end
        3848:
        begin
            RED=8'h60;
            GRN=8'h5D;
            BLU=8'h53;
        end
        3849:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h26;
        end
        3850:
        begin
            RED=8'h2D;
            GRN=8'h2E;
            BLU=8'h26;
        end
        3851:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h28;
        end
        3852:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3853:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3854:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3855:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3856:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3857:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3858:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3859:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3860:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3861:
        begin
            RED=8'h32;
            GRN=8'h33;
            BLU=8'h2B;
        end
        3862:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h28;
        end
        3863:
        begin
            RED=8'h3B;
            GRN=8'h3D;
            BLU=8'h2E;
        end
        3864:
        begin
            RED=8'h6D;
            GRN=8'h6F;
            BLU=8'h62;
        end
        3865:
        begin
            RED=8'hB7;
            GRN=8'hB8;
            BLU=8'hB1;
        end
        3866:
        begin
            RED=8'hF9;
            GRN=8'hFA;
            BLU=8'hF8;
        end
        3867:
        begin
            RED=8'hB7;
            GRN=8'hB2;
            BLU=8'hC0;
        end
        3868:
        begin
            RED=8'h36;
            GRN=8'h21;
            BLU=8'h70;
        end
        3869:
        begin
            RED=8'h36;
            GRN=8'h1C;
            BLU=8'h80;
        end
        3870:
        begin
            RED=8'h35;
            GRN=8'h1B;
            BLU=8'h79;
        end
        3871:
        begin
            RED=8'h36;
            GRN=8'h1C;
            BLU=8'h66;
        end
        3872:
        begin
            RED=8'h69;
            GRN=8'h49;
            BLU=8'h5B;
        end
        3873:
        begin
            RED=8'h9E;
            GRN=8'h7D;
            BLU=8'h84;
        end
        3874:
        begin
            RED=8'h74;
            GRN=8'h52;
            BLU=8'h58;
        end
        3875:
        begin
            RED=8'h80;
            GRN=8'h5E;
            BLU=8'h62;
        end
        3876:
        begin
            RED=8'h7B;
            GRN=8'h5F;
            BLU=8'h73;
        end
        3877:
        begin
            RED=8'h34;
            GRN=8'h20;
            BLU=8'h60;
        end
        3878:
        begin
            RED=8'h34;
            GRN=8'h1C;
            BLU=8'h75;
        end
        3879:
        begin
            RED=8'h37;
            GRN=8'h1C;
            BLU=8'h81;
        end
        3880:
        begin
            RED=8'h38;
            GRN=8'h1E;
            BLU=8'h81;
        end
        3881:
        begin
            RED=8'h39;
            GRN=8'h1C;
            BLU=8'h7C;
        end
        3882:
        begin
            RED=8'h36;
            GRN=8'h1F;
            BLU=8'h79;
        end
        3883:
        begin
            RED=8'h39;
            GRN=8'h33;
            BLU=8'h6A;
        end
        3884:
        begin
            RED=8'hCF;
            GRN=8'hD8;
            BLU=8'hF3;
        end
        3885:
        begin
            RED=8'hCF;
            GRN=8'hDE;
            BLU=8'hFD;
        end
        3886:
        begin
            RED=8'hD1;
            GRN=8'hDF;
            BLU=8'hFA;
        end
        3887:
        begin
            RED=8'hBD;
            GRN=8'hC2;
            BLU=8'hD2;
        end
        3888:
        begin
            RED=8'hF5;
            GRN=8'hF4;
            BLU=8'hF9;
        end
        3889:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFE;
        end
        3890:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFD;
        end
        3891:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        3892:
        begin
            RED=8'hFB;
            GRN=8'hFB;
            BLU=8'hFB;
        end
        3893:
        begin
            RED=8'hDA;
            GRN=8'hDA;
            BLU=8'hDA;
        end
        3894:
        begin
            RED=8'hF3;
            GRN=8'hF3;
            BLU=8'hF3;
        end
        3895:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        3896:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        3897:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        3898:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        3899:
        begin
            RED=8'hFA;
            GRN=8'hFA;
            BLU=8'hF9;
        end
        3900:
        begin
            RED=8'hE2;
            GRN=8'hE3;
            BLU=8'hE0;
        end
        3901:
        begin
            RED=8'h45;
            GRN=8'h46;
            BLU=8'h42;
        end
        3902:
        begin
            RED=8'h2E;
            GRN=8'h2F;
            BLU=8'h29;
        end
        3903:
        begin
            RED=8'h31;
            GRN=8'h32;
            BLU=8'h2A;
        end
        3904:
        begin
            RED=8'hBA;
            GRN=8'hAF;
            BLU=8'h97;
        end
        3905:
        begin
            RED=8'hBB;
            GRN=8'hB1;
            BLU=8'h99;
        end
        3906:
        begin
            RED=8'hBB;
            GRN=8'hB0;
            BLU=8'h98;
        end
        3907:
        begin
            RED=8'hBB;
            GRN=8'hB1;
            BLU=8'h98;
        end
        3908:
        begin
            RED=8'hBA;
            GRN=8'hB1;
            BLU=8'h98;
        end
        3909:
        begin
            RED=8'hB8;
            GRN=8'hB2;
            BLU=8'h98;
        end
        3910:
        begin
            RED=8'hB8;
            GRN=8'hB1;
            BLU=8'h98;
        end
        3911:
        begin
            RED=8'hB7;
            GRN=8'hB0;
            BLU=8'h9A;
        end
        3912:
        begin
            RED=8'hB3;
            GRN=8'hAB;
            BLU=8'h98;
        end
        3913:
        begin
            RED=8'h38;
            GRN=8'h36;
            BLU=8'h2A;
        end
        3914:
        begin
            RED=8'h29;
            GRN=8'h2A;
            BLU=8'h22;
        end
        3915:
        begin
            RED=8'h2D;
            GRN=8'h2E;
            BLU=8'h26;
        end
        3916:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3917:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3918:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3919:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3920:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3921:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3922:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3923:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3924:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h28;
        end
        3925:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3926:
        begin
            RED=8'h31;
            GRN=8'h32;
            BLU=8'h2A;
        end
        3927:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h2B;
        end
        3928:
        begin
            RED=8'h36;
            GRN=8'h36;
            BLU=8'h32;
        end
        3929:
        begin
            RED=8'hE8;
            GRN=8'hE8;
            BLU=8'hE7;
        end
        3930:
        begin
            RED=8'hF9;
            GRN=8'hF9;
            BLU=8'hFB;
        end
        3931:
        begin
            RED=8'hB5;
            GRN=8'hAE;
            BLU=8'hC4;
        end
        3932:
        begin
            RED=8'h37;
            GRN=8'h20;
            BLU=8'h79;
        end
        3933:
        begin
            RED=8'h34;
            GRN=8'h1B;
            BLU=8'h7A;
        end
        3934:
        begin
            RED=8'h38;
            GRN=8'h1E;
            BLU=8'h7C;
        end
        3935:
        begin
            RED=8'h39;
            GRN=8'h1D;
            BLU=8'h7C;
        end
        3936:
        begin
            RED=8'h2F;
            GRN=8'h15;
            BLU=8'h63;
        end
        3937:
        begin
            RED=8'h36;
            GRN=8'h1C;
            BLU=8'h6B;
        end
        3938:
        begin
            RED=8'h36;
            GRN=8'h1C;
            BLU=8'h6B;
        end
        3939:
        begin
            RED=8'h33;
            GRN=8'h1A;
            BLU=8'h62;
        end
        3940:
        begin
            RED=8'h35;
            GRN=8'h1C;
            BLU=8'h69;
        end
        3941:
        begin
            RED=8'h36;
            GRN=8'h1D;
            BLU=8'h78;
        end
        3942:
        begin
            RED=8'h35;
            GRN=8'h1D;
            BLU=8'h74;
        end
        3943:
        begin
            RED=8'h36;
            GRN=8'h1D;
            BLU=8'h79;
        end
        3944:
        begin
            RED=8'h38;
            GRN=8'h1D;
            BLU=8'h83;
        end
        3945:
        begin
            RED=8'h37;
            GRN=8'h1C;
            BLU=8'h7F;
        end
        3946:
        begin
            RED=8'h35;
            GRN=8'h20;
            BLU=8'h76;
        end
        3947:
        begin
            RED=8'h62;
            GRN=8'h5E;
            BLU=8'h8E;
        end
        3948:
        begin
            RED=8'hD2;
            GRN=8'hDE;
            BLU=8'hF6;
        end
        3949:
        begin
            RED=8'hCF;
            GRN=8'hDF;
            BLU=8'hFD;
        end
        3950:
        begin
            RED=8'hD2;
            GRN=8'hE0;
            BLU=8'hFA;
        end
        3951:
        begin
            RED=8'hB2;
            GRN=8'hB7;
            BLU=8'hC4;
        end
        3952:
        begin
            RED=8'hFB;
            GRN=8'hFA;
            BLU=8'hFE;
        end
        3953:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFD;
        end
        3954:
        begin
            RED=8'hFC;
            GRN=8'hFD;
            BLU=8'hFC;
        end
        3955:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        3956:
        begin
            RED=8'hFA;
            GRN=8'hFA;
            BLU=8'hFA;
        end
        3957:
        begin
            RED=8'hD7;
            GRN=8'hD7;
            BLU=8'hD7;
        end
        3958:
        begin
            RED=8'hF5;
            GRN=8'hF5;
            BLU=8'hF5;
        end
        3959:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        3960:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        3961:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        3962:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        3963:
        begin
            RED=8'hFB;
            GRN=8'hFB;
            BLU=8'hFC;
        end
        3964:
        begin
            RED=8'hF8;
            GRN=8'hF8;
            BLU=8'hF8;
        end
        3965:
        begin
            RED=8'hD4;
            GRN=8'hD4;
            BLU=8'hD1;
        end
        3966:
        begin
            RED=8'h34;
            GRN=8'h35;
            BLU=8'h2F;
        end
        3967:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h2A;
        end
        3968:
        begin
            RED=8'hBB;
            GRN=8'hB1;
            BLU=8'h96;
        end
        3969:
        begin
            RED=8'hBB;
            GRN=8'hB1;
            BLU=8'h96;
        end
        3970:
        begin
            RED=8'hBB;
            GRN=8'hB1;
            BLU=8'h96;
        end
        3971:
        begin
            RED=8'hBB;
            GRN=8'hB1;
            BLU=8'h96;
        end
        3972:
        begin
            RED=8'hBA;
            GRN=8'hB1;
            BLU=8'h96;
        end
        3973:
        begin
            RED=8'hB8;
            GRN=8'hB3;
            BLU=8'h94;
        end
        3974:
        begin
            RED=8'hB8;
            GRN=8'hB2;
            BLU=8'h95;
        end
        3975:
        begin
            RED=8'hB8;
            GRN=8'hB2;
            BLU=8'h97;
        end
        3976:
        begin
            RED=8'hB4;
            GRN=8'hAC;
            BLU=8'h94;
        end
        3977:
        begin
            RED=8'h3D;
            GRN=8'h3B;
            BLU=8'h2E;
        end
        3978:
        begin
            RED=8'h2B;
            GRN=8'h2C;
            BLU=8'h24;
        end
        3979:
        begin
            RED=8'h27;
            GRN=8'h28;
            BLU=8'h20;
        end
        3980:
        begin
            RED=8'h2A;
            GRN=8'h2B;
            BLU=8'h23;
        end
        3981:
        begin
            RED=8'h2E;
            GRN=8'h2F;
            BLU=8'h27;
        end
        3982:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3983:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3984:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3985:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3986:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3987:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3988:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3989:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        3990:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h2A;
        end
        3991:
        begin
            RED=8'h30;
            GRN=8'h30;
            BLU=8'h2D;
        end
        3992:
        begin
            RED=8'h48;
            GRN=8'h48;
            BLU=8'h46;
        end
        3993:
        begin
            RED=8'hF7;
            GRN=8'hF7;
            BLU=8'hF5;
        end
        3994:
        begin
            RED=8'hFB;
            GRN=8'hFB;
            BLU=8'hFA;
        end
        3995:
        begin
            RED=8'hE0;
            GRN=8'hDC;
            BLU=8'hE5;
        end
        3996:
        begin
            RED=8'h38;
            GRN=8'h25;
            BLU=8'h6B;
        end
        3997:
        begin
            RED=8'h34;
            GRN=8'h1D;
            BLU=8'h73;
        end
        3998:
        begin
            RED=8'h30;
            GRN=8'h17;
            BLU=8'h6F;
        end
        3999:
        begin
            RED=8'h2E;
            GRN=8'h14;
            BLU=8'h66;
        end
        4000:
        begin
            RED=8'h2E;
            GRN=8'h19;
            BLU=8'h66;
        end
        4001:
        begin
            RED=8'h34;
            GRN=8'h1F;
            BLU=8'h76;
        end
        4002:
        begin
            RED=8'h35;
            GRN=8'h1F;
            BLU=8'h78;
        end
        4003:
        begin
            RED=8'h2C;
            GRN=8'h18;
            BLU=8'h67;
        end
        4004:
        begin
            RED=8'h2E;
            GRN=8'h19;
            BLU=8'h66;
        end
        4005:
        begin
            RED=8'h32;
            GRN=8'h1A;
            BLU=8'h72;
        end
        4006:
        begin
            RED=8'h32;
            GRN=8'h1B;
            BLU=8'h6E;
        end
        4007:
        begin
            RED=8'h35;
            GRN=8'h1D;
            BLU=8'h72;
        end
        4008:
        begin
            RED=8'h37;
            GRN=8'h1E;
            BLU=8'h79;
        end
        4009:
        begin
            RED=8'h37;
            GRN=8'h1D;
            BLU=8'h7E;
        end
        4010:
        begin
            RED=8'h32;
            GRN=8'h20;
            BLU=8'h72;
        end
        4011:
        begin
            RED=8'h90;
            GRN=8'h91;
            BLU=8'hBA;
        end
        4012:
        begin
            RED=8'hD1;
            GRN=8'hDF;
            BLU=8'hF3;
        end
        4013:
        begin
            RED=8'hCD;
            GRN=8'hDF;
            BLU=8'hFD;
        end
        4014:
        begin
            RED=8'hCF;
            GRN=8'hDD;
            BLU=8'hF4;
        end
        4015:
        begin
            RED=8'hB8;
            GRN=8'hBE;
            BLU=8'hC9;
        end
        4016:
        begin
            RED=8'hFB;
            GRN=8'hFB;
            BLU=8'hFD;
        end
        4017:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFA;
        end
        4018:
        begin
            RED=8'hFD;
            GRN=8'hFD;
            BLU=8'hFC;
        end
        4019:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        4020:
        begin
            RED=8'hFB;
            GRN=8'hFB;
            BLU=8'hFB;
        end
        4021:
        begin
            RED=8'hC8;
            GRN=8'hC8;
            BLU=8'hC8;
        end
        4022:
        begin
            RED=8'hF9;
            GRN=8'hF9;
            BLU=8'hF9;
        end
        4023:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        4024:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        4025:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        4026:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        4027:
        begin
            RED=8'hFD;
            GRN=8'hFD;
            BLU=8'hFE;
        end
        4028:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFE;
        end
        4029:
        begin
            RED=8'hFA;
            GRN=8'hFA;
            BLU=8'hFA;
        end
        4030:
        begin
            RED=8'hA4;
            GRN=8'hA5;
            BLU=8'hA2;
        end
        4031:
        begin
            RED=8'h2E;
            GRN=8'h2F;
            BLU=8'h2A;
        end
        4032:
        begin
            RED=8'hBA;
            GRN=8'hB4;
            BLU=8'h99;
        end
        4033:
        begin
            RED=8'hB9;
            GRN=8'hB4;
            BLU=8'h99;
        end
        4034:
        begin
            RED=8'hB9;
            GRN=8'hB4;
            BLU=8'h9A;
        end
        4035:
        begin
            RED=8'hB9;
            GRN=8'hB4;
            BLU=8'h9A;
        end
        4036:
        begin
            RED=8'hB9;
            GRN=8'hB5;
            BLU=8'h99;
        end
        4037:
        begin
            RED=8'hB8;
            GRN=8'hB6;
            BLU=8'h97;
        end
        4038:
        begin
            RED=8'hB8;
            GRN=8'hB5;
            BLU=8'h98;
        end
        4039:
        begin
            RED=8'hB7;
            GRN=8'hB5;
            BLU=8'h99;
        end
        4040:
        begin
            RED=8'hB3;
            GRN=8'hAF;
            BLU=8'h97;
        end
        4041:
        begin
            RED=8'h3C;
            GRN=8'h3C;
            BLU=8'h2F;
        end
        4042:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h28;
        end
        4043:
        begin
            RED=8'h2F;
            GRN=8'h30;
            BLU=8'h28;
        end
        4044:
        begin
            RED=8'h2A;
            GRN=8'h2B;
            BLU=8'h23;
        end
        4045:
        begin
            RED=8'h26;
            GRN=8'h28;
            BLU=8'h1F;
        end
        4046:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        4047:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        4048:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        4049:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        4050:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        4051:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        4052:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        4053:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h29;
        end
        4054:
        begin
            RED=8'h30;
            GRN=8'h31;
            BLU=8'h2A;
        end
        4055:
        begin
            RED=8'h2E;
            GRN=8'h2F;
            BLU=8'h2B;
        end
        4056:
        begin
            RED=8'h72;
            GRN=8'h73;
            BLU=8'h6E;
        end
        4057:
        begin
            RED=8'hFC;
            GRN=8'hFD;
            BLU=8'hF7;
        end
        4058:
        begin
            RED=8'hFD;
            GRN=8'hFE;
            BLU=8'hF7;
        end
        4059:
        begin
            RED=8'hF7;
            GRN=8'hF4;
            BLU=8'hF3;
        end
        4060:
        begin
            RED=8'h4E;
            GRN=8'h3B;
            BLU=8'h7A;
        end
        4061:
        begin
            RED=8'h34;
            GRN=8'h1B;
            BLU=8'h7C;
        end
        4062:
        begin
            RED=8'h37;
            GRN=8'h1C;
            BLU=8'h7C;
        end
        4063:
        begin
            RED=8'h32;
            GRN=8'h1A;
            BLU=8'h63;
        end
        4064:
        begin
            RED=8'h35;
            GRN=8'h1D;
            BLU=8'h6A;
        end
        4065:
        begin
            RED=8'h38;
            GRN=8'h1E;
            BLU=8'h7B;
        end
        4066:
        begin
            RED=8'h38;
            GRN=8'h1E;
            BLU=8'h7E;
        end
        4067:
        begin
            RED=8'h32;
            GRN=8'h1A;
            BLU=8'h6E;
        end
        4068:
        begin
            RED=8'h35;
            GRN=8'h1D;
            BLU=8'h69;
        end
        4069:
        begin
            RED=8'h33;
            GRN=8'h1B;
            BLU=8'h72;
        end
        4070:
        begin
            RED=8'h34;
            GRN=8'h1A;
            BLU=8'h7C;
        end
        4071:
        begin
            RED=8'h35;
            GRN=8'h1A;
            BLU=8'h7F;
        end
        4072:
        begin
            RED=8'h37;
            GRN=8'h1D;
            BLU=8'h7D;
        end
        4073:
        begin
            RED=8'h36;
            GRN=8'h1E;
            BLU=8'h7E;
        end
        4074:
        begin
            RED=8'h32;
            GRN=8'h22;
            BLU=8'h71;
        end
        4075:
        begin
            RED=8'hA7;
            GRN=8'hA9;
            BLU=8'hCE;
        end
        4076:
        begin
            RED=8'hD0;
            GRN=8'hE0;
            BLU=8'hF2;
        end
        4077:
        begin
            RED=8'hCD;
            GRN=8'hE1;
            BLU=8'hFE;
        end
        4078:
        begin
            RED=8'hCE;
            GRN=8'hDC;
            BLU=8'hF2;
        end
        4079:
        begin
            RED=8'hCE;
            GRN=8'hD3;
            BLU=8'hDA;
        end
        4080:
        begin
            RED=8'hFB;
            GRN=8'hFB;
            BLU=8'hFC;
        end
        4081:
        begin
            RED=8'hFC;
            GRN=8'hFD;
            BLU=8'hF9;
        end
        4082:
        begin
            RED=8'hFD;
            GRN=8'hFD;
            BLU=8'hFC;
        end
        4083:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        4084:
        begin
            RED=8'hFA;
            GRN=8'hFA;
            BLU=8'hFA;
        end
        4085:
        begin
            RED=8'hC9;
            GRN=8'hC9;
            BLU=8'hC9;
        end
        4086:
        begin
            RED=8'hF9;
            GRN=8'hF9;
            BLU=8'hF9;
        end
        4087:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        4088:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        4089:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        4090:
        begin
            RED=8'hFC;
            GRN=8'hFC;
            BLU=8'hFC;
        end
        4091:
        begin
            RED=8'hFD;
            GRN=8'hFC;
            BLU=8'hFE;
        end
        4092:
        begin
            RED=8'hFC;
            GRN=8'hFB;
            BLU=8'hFF;
        end
        4093:
        begin
            RED=8'hFB;
            GRN=8'hFB;
            BLU=8'hFD;
        end
        4094:
        begin
            RED=8'hF2;
            GRN=8'hF2;
            BLU=8'hF1;
        end
        4095:
        begin
            RED=8'h5E;
            GRN=8'h5E;
            BLU=8'h5B;
        end
        default:
        begin
            RED=8'h00;
            GRN=8'h00;
            BLU=8'h00;
        end
    endcase
endmodule
